module debug_log(
	input clock, reset,
	input[7:0] data,
	output TXD
);


endmodule
