// Generator : SpinalHDL v1.4.3    git head : adf552d8f500e7419fff395b7049228e4bc5de26
// Component : TopLevel
// Git hash  : 2ed321ce8dc266500e84f5d75b457f0baa0e827d


`define machine_enumDefinition_defaultEncoding_type [2:0]
`define machine_enumDefinition_defaultEncoding_machine_BOOT 3'b000
`define machine_enumDefinition_defaultEncoding_machine_idle 3'b001
`define machine_enumDefinition_defaultEncoding_machine_init 3'b010
`define machine_enumDefinition_defaultEncoding_machine_tx 3'b011
`define machine_enumDefinition_defaultEncoding_machine_rx 3'b100
`define machine_enumDefinition_defaultEncoding_machine_ack 3'b101

`define UartParityType_defaultEncoding_type [1:0]
`define UartParityType_defaultEncoding_NONE 2'b00
`define UartParityType_defaultEncoding_EVEN 2'b01
`define UartParityType_defaultEncoding_ODD 2'b10

`define UartStopType_defaultEncoding_type [0:0]
`define UartStopType_defaultEncoding_ONE 1'b0
`define UartStopType_defaultEncoding_TWO 1'b1

`define machine_enumDefinition_1_defaultEncoding_type [3:0]
`define machine_enumDefinition_1_defaultEncoding_machine_BOOT 4'b0000
`define machine_enumDefinition_1_defaultEncoding_machine_idle 4'b0001
`define machine_enumDefinition_1_defaultEncoding_machine_k6 4'b0010
`define machine_enumDefinition_1_defaultEncoding_machine_k5 4'b0011
`define machine_enumDefinition_1_defaultEncoding_machine_k4 4'b0100
`define machine_enumDefinition_1_defaultEncoding_machine_k3 4'b0101
`define machine_enumDefinition_1_defaultEncoding_machine_k2 4'b0110
`define machine_enumDefinition_1_defaultEncoding_machine_k1 4'b0111
`define machine_enumDefinition_1_defaultEncoding_machine_reserved 4'b1000
`define machine_enumDefinition_1_defaultEncoding_machine_special 4'b1001

`define UartCtrlTxState_defaultEncoding_type [2:0]
`define UartCtrlTxState_defaultEncoding_IDLE 3'b000
`define UartCtrlTxState_defaultEncoding_START 3'b001
`define UartCtrlTxState_defaultEncoding_DATA 3'b010
`define UartCtrlTxState_defaultEncoding_PARITY 3'b011
`define UartCtrlTxState_defaultEncoding_STOP 3'b100

`define UartCtrlRxState_defaultEncoding_type [2:0]
`define UartCtrlRxState_defaultEncoding_IDLE 3'b000
`define UartCtrlRxState_defaultEncoding_START 3'b001
`define UartCtrlRxState_defaultEncoding_DATA 3'b010
`define UartCtrlRxState_defaultEncoding_PARITY 3'b011
`define UartCtrlRxState_defaultEncoding_STOP 3'b100


module TopLevel (
  input               KEY_Fn,
  input               CLK_50,
  input      [20:0]   COL,
  output     [5:0]    LED_A,
  output     [5:0]    ROW,
  output     [34:0]   LED_K,
  output              TXD,
  output              LED_R6,
   inout              PS2_CLK,
   inout              PS2_DAT
);
  wire                _zz_3;
  wire                _zz_4;
  wire                _zz_5;
  wire                _zz_6;
  wire                rstCtrl_io_globalReset;
  wire       [5:0]    core_led_row_export;
  wire       [34:0]   core_led_col_export;
  wire                core_send_to_host_valid;
  wire       [7:0]    core_send_to_host_payload;
  wire                core_receive_from_host_ready;
  wire                core_locked_export;
  wire                bufferCC_2_io_dataOut;
  wire       [5:0]    clk50Area_keyMatrix_ROW;
  wire                clk50Area_keyMatrix_scanIdx_valid;
  wire       [7:0]    clk50Area_keyMatrix_scanIdx_payload;
  wire       [205:0]  clk50Area_keyMatrix_keyBits;
  wire                clk50Area_ps2_receiveFromHost_valid;
  wire       [7:0]    clk50Area_ps2_receiveFromHost_payload;
  wire                clk50Area_ps2_sendToHost_ready;
  wire                clk50Area_hid_TXD;
  reg                 _zz_1;
  wire                _zz_2;

  ResetController rstCtrl (
    .io_clock            (CLK_50                  ), //i
    .io_externalReset    (_zz_3                   ), //i
    .io_globalReset      (rstCtrl_io_globalReset  )  //o
  );
  TPK core (
    .clk_clk                      (CLK_50                                      ), //i
    .reset_reset_n                (_zz_4                                       ), //i
    .led_row_export               (core_led_row_export[5:0]                    ), //o
    .led_col_export               (core_led_col_export[34:0]                   ), //o
    .scan_idx_valid               (clk50Area_keyMatrix_scanIdx_valid           ), //i
    .scan_idx_payload             (clk50Area_keyMatrix_scanIdx_payload[7:0]    ), //i
    .send_to_host_valid           (core_send_to_host_valid                     ), //o
    .send_to_host_ready           (clk50Area_ps2_sendToHost_ready              ), //i
    .send_to_host_payload         (core_send_to_host_payload[7:0]              ), //o
    .receive_from_host_valid      (clk50Area_ps2_receiveFromHost_valid         ), //i
    .receive_from_host_ready      (core_receive_from_host_ready                ), //o
    .receive_from_host_payload    (clk50Area_ps2_receiveFromHost_payload[7:0]  ), //i
    .locked_export                (core_locked_export                          )  //o
  );
  BufferCC_1 bufferCC_2 (
    .io_dataIn     (_zz_5                  ), //i
    .io_dataOut    (bufferCC_2_io_dataOut  ), //o
    .CLK_50        (CLK_50                 ), //i
    ._zz_1         (_zz_2                  )  //i
  );
  KeyMatrix clk50Area_keyMatrix (
    .enabled            (_zz_6                                     ), //i
    .COL                (COL[20:0]                                 ), //i
    .ROW                (clk50Area_keyMatrix_ROW[5:0]              ), //o
    .scanIdx_valid      (clk50Area_keyMatrix_scanIdx_valid         ), //o
    .scanIdx_payload    (clk50Area_keyMatrix_scanIdx_payload[7:0]  ), //o
    .keyBits            (clk50Area_keyMatrix_keyBits[205:0]        ), //o
    ._zz_1              (_zz_1                                     ), //i
    .CLK_50             (CLK_50                                    )  //i
  );
  PS2Device clk50Area_ps2 (
    .PS2_CLK                    (PS2_CLK                                     ), //~
    .PS2_DAT                    (PS2_DAT                                     ), //~
    .receiveFromHost_valid      (clk50Area_ps2_receiveFromHost_valid         ), //o
    .receiveFromHost_payload    (clk50Area_ps2_receiveFromHost_payload[7:0]  ), //o
    .sendToHost_valid           (core_send_to_host_valid                     ), //i
    .sendToHost_ready           (clk50Area_ps2_sendToHost_ready              ), //o
    .sendToHost_payload         (core_send_to_host_payload[7:0]              ), //i
    ._zz_3                      (_zz_1                                       ), //i
    .CLK_50                     (CLK_50                                      )  //i
  );
  HID clk50Area_hid (
    .TXD                (clk50Area_hid_TXD                         ), //o
    .scanIdx_valid      (clk50Area_keyMatrix_scanIdx_valid         ), //i
    .scanIdx_payload    (clk50Area_keyMatrix_scanIdx_payload[7:0]  ), //i
    .keyBits            (clk50Area_keyMatrix_keyBits[205:0]        ), //i
    .CLK_50             (CLK_50                                    ), //i
    ._zz_104            (_zz_1                                     )  //i
  );
  assign _zz_3 = (! KEY_Fn);
  always @ (*) begin
    _zz_1 = 1'b0;
    _zz_1 = bufferCC_2_io_dataOut;
  end

  assign _zz_4 = (! _zz_1);
  assign _zz_2 = (rstCtrl_io_globalReset || (! core_locked_export));
  assign _zz_5 = 1'b0;
  assign LED_A = core_led_row_export;
  assign LED_K = core_led_col_export;
  assign LED_R6 = 1'b1;
  assign ROW = clk50Area_keyMatrix_ROW;
  assign _zz_6 = 1'b1;
  assign TXD = clk50Area_hid_TXD;

endmodule

module HID (
  output              TXD,
  input               scanIdx_valid,
  input      [7:0]    scanIdx_payload,
  input      [205:0]  keyBits,
  input               CLK_50,
  input               _zz_104
);
  wire       [2:0]    _zz_105;
  wire       `UartStopType_defaultEncoding_type _zz_106;
  wire       `UartParityType_defaultEncoding_type _zz_107;
  wire       [19:0]   _zz_108;
  wire                _zz_109;
  reg        [7:0]    _zz_110;
  wire                _zz_111;
  wire                _zz_112;
  wire                _zz_113;
  reg        [7:0]    _zz_114;
  wire                uartCtrl_1_io_write_ready;
  wire                uartCtrl_1_io_read_valid;
  wire       [7:0]    uartCtrl_1_io_read_payload;
  wire                uartCtrl_1_io_uart_txd;
  wire                uartCtrl_1_io_readError;
  wire                uartCtrl_1_io_readBreak;
  wire       [0:0]    _zz_115;
  wire       [0:0]    _zz_116;
  wire       [0:0]    _zz_117;
  wire       [0:0]    _zz_118;
  wire       [0:0]    _zz_119;
  wire       [0:0]    _zz_120;
  wire       [0:0]    _zz_121;
  wire       [0:0]    _zz_122;
  wire       [0:0]    _zz_123;
  wire       [0:0]    _zz_124;
  wire       [0:0]    _zz_125;
  wire       [0:0]    _zz_126;
  wire       [0:0]    _zz_127;
  wire       [0:0]    _zz_128;
  wire       [0:0]    _zz_129;
  wire       [0:0]    _zz_130;
  wire       [0:0]    _zz_131;
  wire       [0:0]    _zz_132;
  wire       [0:0]    _zz_133;
  wire       [0:0]    _zz_134;
  wire       [0:0]    _zz_135;
  wire       [0:0]    _zz_136;
  wire       [0:0]    _zz_137;
  wire       [0:0]    _zz_138;
  wire       [0:0]    _zz_139;
  wire       [0:0]    _zz_140;
  wire       [0:0]    _zz_141;
  wire       [0:0]    _zz_142;
  wire       [0:0]    _zz_143;
  wire       [0:0]    _zz_144;
  wire       [0:0]    _zz_145;
  wire       [0:0]    _zz_146;
  wire       [0:0]    _zz_147;
  wire       [0:0]    _zz_148;
  wire       [0:0]    _zz_149;
  wire       [0:0]    _zz_150;
  wire       [0:0]    _zz_151;
  wire       [0:0]    _zz_152;
  wire       [0:0]    _zz_153;
  wire       [0:0]    _zz_154;
  wire       [0:0]    _zz_155;
  wire       [0:0]    _zz_156;
  wire       [0:0]    _zz_157;
  wire       [0:0]    _zz_158;
  wire       [0:0]    _zz_159;
  wire       [0:0]    _zz_160;
  wire       [0:0]    _zz_161;
  wire       [0:0]    _zz_162;
  wire       [0:0]    _zz_163;
  wire       [0:0]    _zz_164;
  wire       [0:0]    _zz_165;
  wire       [0:0]    _zz_166;
  wire       [0:0]    _zz_167;
  wire       [0:0]    _zz_168;
  wire       [0:0]    _zz_169;
  wire       [0:0]    _zz_170;
  wire       [0:0]    _zz_171;
  wire       [0:0]    _zz_172;
  wire       [0:0]    _zz_173;
  wire       [0:0]    _zz_174;
  wire       [0:0]    _zz_175;
  wire       [0:0]    _zz_176;
  wire       [0:0]    _zz_177;
  wire       [0:0]    _zz_178;
  wire       [0:0]    _zz_179;
  wire       [0:0]    _zz_180;
  wire       [0:0]    _zz_181;
  wire       [0:0]    _zz_182;
  wire       [0:0]    _zz_183;
  wire       [0:0]    _zz_184;
  wire       [0:0]    _zz_185;
  wire       [0:0]    _zz_186;
  wire       [0:0]    _zz_187;
  wire       [0:0]    _zz_188;
  wire       [0:0]    _zz_189;
  wire       [0:0]    _zz_190;
  wire       [0:0]    _zz_191;
  wire       [0:0]    _zz_192;
  wire       [0:0]    _zz_193;
  wire       [0:0]    _zz_194;
  wire       [0:0]    _zz_195;
  wire       [0:0]    _zz_196;
  wire       [0:0]    _zz_197;
  wire       [0:0]    _zz_198;
  wire       [0:0]    _zz_199;
  wire       [0:0]    _zz_200;
  wire       [0:0]    _zz_201;
  wire       [0:0]    _zz_202;
  wire       [0:0]    _zz_203;
  wire       [0:0]    _zz_204;
  wire       [0:0]    _zz_205;
  wire       [0:0]    _zz_206;
  wire       [0:0]    _zz_207;
  wire       [0:0]    _zz_208;
  wire       [0:0]    _zz_209;
  wire       [0:0]    _zz_210;
  wire       [0:0]    _zz_211;
  wire       [0:0]    _zz_212;
  wire       [0:0]    _zz_213;
  wire       [0:0]    _zz_214;
  wire       [0:0]    _zz_215;
  wire       [0:0]    _zz_216;
  wire       [0:0]    _zz_217;
  wire       [0:0]    _zz_218;
  wire       [0:0]    _zz_219;
  wire       [0:0]    _zz_220;
  wire       [0:0]    _zz_221;
  wire       [0:0]    _zz_222;
  wire       [0:0]    _zz_223;
  wire       [0:0]    _zz_224;
  wire       [0:0]    _zz_225;
  wire       [0:0]    _zz_226;
  wire       [0:0]    _zz_227;
  wire       [0:0]    _zz_228;
  wire       [0:0]    _zz_229;
  wire       [0:0]    _zz_230;
  wire       [0:0]    _zz_231;
  wire       [0:0]    _zz_232;
  wire       [0:0]    _zz_233;
  wire       [0:0]    _zz_234;
  wire       [0:0]    _zz_235;
  wire       [0:0]    _zz_236;
  wire       [0:0]    _zz_237;
  wire       [0:0]    _zz_238;
  wire       [0:0]    _zz_239;
  wire       [0:0]    _zz_240;
  wire       [0:0]    _zz_241;
  wire       [0:0]    _zz_242;
  wire       [0:0]    _zz_243;
  wire       [0:0]    _zz_244;
  wire       [0:0]    _zz_245;
  wire       [0:0]    _zz_246;
  wire       [0:0]    _zz_247;
  wire       [0:0]    _zz_248;
  wire       [0:0]    _zz_249;
  wire       [0:0]    _zz_250;
  wire       [0:0]    _zz_251;
  wire       [0:0]    _zz_252;
  wire       [0:0]    _zz_253;
  wire       [0:0]    _zz_254;
  wire       [0:0]    _zz_255;
  wire       [0:0]    _zz_256;
  wire       [0:0]    _zz_257;
  wire       [0:0]    _zz_258;
  wire       [0:0]    _zz_259;
  wire       [0:0]    _zz_260;
  wire       [0:0]    _zz_261;
  wire       [0:0]    _zz_262;
  wire       [0:0]    _zz_263;
  wire       [0:0]    _zz_264;
  wire       [0:0]    _zz_265;
  wire       [0:0]    _zz_266;
  wire       [0:0]    _zz_267;
  wire       [0:0]    _zz_268;
  wire       [0:0]    _zz_269;
  wire       [0:0]    _zz_270;
  wire       [0:0]    _zz_271;
  wire       [0:0]    _zz_272;
  wire       [0:0]    _zz_273;
  wire       [0:0]    _zz_274;
  wire       [0:0]    _zz_275;
  wire       [0:0]    _zz_276;
  wire       [0:0]    _zz_277;
  wire       [0:0]    _zz_278;
  wire       [0:0]    _zz_279;
  wire       [0:0]    _zz_280;
  wire       [0:0]    _zz_281;
  wire       [0:0]    _zz_282;
  wire       [0:0]    _zz_283;
  wire       [0:0]    _zz_284;
  wire       [0:0]    _zz_285;
  wire       [0:0]    _zz_286;
  wire       [0:0]    _zz_287;
  wire       [0:0]    _zz_288;
  wire       [0:0]    _zz_289;
  wire       [0:0]    _zz_290;
  wire       [0:0]    _zz_291;
  wire       [0:0]    _zz_292;
  wire       [0:0]    _zz_293;
  wire       [0:0]    _zz_294;
  wire       [0:0]    _zz_295;
  wire       [0:0]    _zz_296;
  wire       [0:0]    _zz_297;
  wire       [0:0]    _zz_298;
  wire       [0:0]    _zz_299;
  wire       [0:0]    _zz_300;
  wire       [0:0]    _zz_301;
  wire       [0:0]    _zz_302;
  wire       [0:0]    _zz_303;
  wire       [0:0]    _zz_304;
  wire       [0:0]    _zz_305;
  wire       [0:0]    _zz_306;
  wire       [0:0]    _zz_307;
  wire       [0:0]    _zz_308;
  wire       [0:0]    _zz_309;
  wire       [0:0]    _zz_310;
  wire       [0:0]    _zz_311;
  wire       [0:0]    _zz_312;
  wire       [0:0]    _zz_313;
  wire       [0:0]    _zz_314;
  wire       [0:0]    _zz_315;
  wire       [0:0]    _zz_316;
  wire       [0:0]    _zz_317;
  wire       [0:0]    _zz_318;
  wire       [0:0]    _zz_319;
  wire       [0:0]    _zz_320;
  wire                _zz_321;
  wire                keyStatus_0_valid;
  wire                keyStatus_0_payload;
  wire                keyStatus_1_valid;
  wire                keyStatus_1_payload;
  wire                keyStatus_2_valid;
  wire                keyStatus_2_payload;
  wire                keyStatus_3_valid;
  wire                keyStatus_3_payload;
  wire                keyStatus_4_valid;
  wire                keyStatus_4_payload;
  wire                keyStatus_5_valid;
  wire                keyStatus_5_payload;
  wire                keyStatus_6_valid;
  wire                keyStatus_6_payload;
  wire                keyStatus_7_valid;
  wire                keyStatus_7_payload;
  wire                keyStatus_8_valid;
  wire                keyStatus_8_payload;
  wire                keyStatus_9_valid;
  wire                keyStatus_9_payload;
  wire                keyStatus_10_valid;
  wire                keyStatus_10_payload;
  wire                keyStatus_11_valid;
  wire                keyStatus_11_payload;
  wire                keyStatus_12_valid;
  wire                keyStatus_12_payload;
  wire                keyStatus_13_valid;
  wire                keyStatus_13_payload;
  wire                keyStatus_14_valid;
  wire                keyStatus_14_payload;
  wire                keyStatus_15_valid;
  wire                keyStatus_15_payload;
  wire                keyStatus_16_valid;
  wire                keyStatus_16_payload;
  wire                keyStatus_17_valid;
  wire                keyStatus_17_payload;
  wire                keyStatus_18_valid;
  wire                keyStatus_18_payload;
  wire                keyStatus_19_valid;
  wire                keyStatus_19_payload;
  wire                keyStatus_20_valid;
  wire                keyStatus_20_payload;
  wire                keyStatus_21_valid;
  wire                keyStatus_21_payload;
  wire                keyStatus_22_valid;
  wire                keyStatus_22_payload;
  wire                keyStatus_23_valid;
  wire                keyStatus_23_payload;
  wire                keyStatus_24_valid;
  wire                keyStatus_24_payload;
  wire                keyStatus_25_valid;
  wire                keyStatus_25_payload;
  wire                keyStatus_26_valid;
  wire                keyStatus_26_payload;
  wire                keyStatus_27_valid;
  wire                keyStatus_27_payload;
  wire                keyStatus_28_valid;
  wire                keyStatus_28_payload;
  wire                keyStatus_29_valid;
  wire                keyStatus_29_payload;
  wire                keyStatus_30_valid;
  wire                keyStatus_30_payload;
  wire                keyStatus_31_valid;
  wire                keyStatus_31_payload;
  wire                keyStatus_32_valid;
  wire                keyStatus_32_payload;
  wire                keyStatus_33_valid;
  wire                keyStatus_33_payload;
  wire                keyStatus_34_valid;
  wire                keyStatus_34_payload;
  wire                keyStatus_35_valid;
  wire                keyStatus_35_payload;
  wire                keyStatus_36_valid;
  wire                keyStatus_36_payload;
  wire                keyStatus_37_valid;
  wire                keyStatus_37_payload;
  wire                keyStatus_38_valid;
  wire                keyStatus_38_payload;
  wire                keyStatus_39_valid;
  wire                keyStatus_39_payload;
  wire                keyStatus_40_valid;
  wire                keyStatus_40_payload;
  wire                keyStatus_41_valid;
  wire                keyStatus_41_payload;
  wire                keyStatus_42_valid;
  wire                keyStatus_42_payload;
  wire                keyStatus_43_valid;
  wire                keyStatus_43_payload;
  wire                keyStatus_44_valid;
  wire                keyStatus_44_payload;
  wire                keyStatus_45_valid;
  wire                keyStatus_45_payload;
  wire                keyStatus_46_valid;
  wire                keyStatus_46_payload;
  wire                keyStatus_47_valid;
  wire                keyStatus_47_payload;
  wire                keyStatus_48_valid;
  wire                keyStatus_48_payload;
  wire                keyStatus_49_valid;
  wire                keyStatus_49_payload;
  wire                keyStatus_50_valid;
  wire                keyStatus_50_payload;
  wire                keyStatus_51_valid;
  wire                keyStatus_51_payload;
  wire                keyStatus_52_valid;
  wire                keyStatus_52_payload;
  wire                keyStatus_53_valid;
  wire                keyStatus_53_payload;
  wire                keyStatus_54_valid;
  wire                keyStatus_54_payload;
  wire                keyStatus_55_valid;
  wire                keyStatus_55_payload;
  wire                keyStatus_56_valid;
  wire                keyStatus_56_payload;
  wire                keyStatus_57_valid;
  wire                keyStatus_57_payload;
  wire                keyStatus_58_valid;
  wire                keyStatus_58_payload;
  wire                keyStatus_59_valid;
  wire                keyStatus_59_payload;
  wire                keyStatus_60_valid;
  wire                keyStatus_60_payload;
  wire                keyStatus_61_valid;
  wire                keyStatus_61_payload;
  wire                keyStatus_62_valid;
  wire                keyStatus_62_payload;
  wire                keyStatus_63_valid;
  wire                keyStatus_63_payload;
  wire                keyStatus_64_valid;
  wire                keyStatus_64_payload;
  wire                keyStatus_65_valid;
  wire                keyStatus_65_payload;
  wire                keyStatus_66_valid;
  wire                keyStatus_66_payload;
  wire                keyStatus_67_valid;
  wire                keyStatus_67_payload;
  wire                keyStatus_68_valid;
  wire                keyStatus_68_payload;
  wire                keyStatus_69_valid;
  wire                keyStatus_69_payload;
  wire                keyStatus_70_valid;
  wire                keyStatus_70_payload;
  wire                keyStatus_71_valid;
  wire                keyStatus_71_payload;
  wire                keyStatus_72_valid;
  wire                keyStatus_72_payload;
  wire                keyStatus_73_valid;
  wire                keyStatus_73_payload;
  wire                keyStatus_74_valid;
  wire                keyStatus_74_payload;
  wire                keyStatus_75_valid;
  wire                keyStatus_75_payload;
  wire                keyStatus_76_valid;
  wire                keyStatus_76_payload;
  wire                keyStatus_77_valid;
  wire                keyStatus_77_payload;
  wire                keyStatus_78_valid;
  wire                keyStatus_78_payload;
  wire                keyStatus_79_valid;
  wire                keyStatus_79_payload;
  wire                keyStatus_80_valid;
  wire                keyStatus_80_payload;
  wire                keyStatus_81_valid;
  wire                keyStatus_81_payload;
  wire                keyStatus_82_valid;
  wire                keyStatus_82_payload;
  wire                keyStatus_83_valid;
  wire                keyStatus_83_payload;
  wire                keyStatus_84_valid;
  wire                keyStatus_84_payload;
  wire                keyStatus_85_valid;
  wire                keyStatus_85_payload;
  wire                keyStatus_86_valid;
  wire                keyStatus_86_payload;
  wire                keyStatus_87_valid;
  wire                keyStatus_87_payload;
  wire                keyStatus_88_valid;
  wire                keyStatus_88_payload;
  wire                keyStatus_89_valid;
  wire                keyStatus_89_payload;
  wire                keyStatus_90_valid;
  wire                keyStatus_90_payload;
  wire                keyStatus_91_valid;
  wire                keyStatus_91_payload;
  wire                keyStatus_92_valid;
  wire                keyStatus_92_payload;
  wire                keyStatus_93_valid;
  wire                keyStatus_93_payload;
  wire                keyStatus_94_valid;
  wire                keyStatus_94_payload;
  wire                keyStatus_95_valid;
  wire                keyStatus_95_payload;
  wire                keyStatus_96_valid;
  wire                keyStatus_96_payload;
  wire                keyStatus_97_valid;
  wire                keyStatus_97_payload;
  wire                keyStatus_98_valid;
  wire                keyStatus_98_payload;
  wire                keyStatus_99_valid;
  wire                keyStatus_99_payload;
  wire                keyStatus_100_valid;
  wire                keyStatus_100_payload;
  wire                keyStatus_101_valid;
  wire                keyStatus_101_payload;
  wire                keyStatus_102_valid;
  wire                keyStatus_102_payload;
  wire       [1:0]    _zz_1;
  wire       [1:0]    _zz_2;
  wire       [1:0]    _zz_3;
  wire       [1:0]    _zz_4;
  wire       [1:0]    _zz_5;
  wire       [1:0]    _zz_6;
  wire       [1:0]    _zz_7;
  wire       [1:0]    _zz_8;
  wire       [1:0]    _zz_9;
  wire       [1:0]    _zz_10;
  wire       [1:0]    _zz_11;
  wire       [1:0]    _zz_12;
  wire       [1:0]    _zz_13;
  wire       [1:0]    _zz_14;
  wire       [1:0]    _zz_15;
  wire       [1:0]    _zz_16;
  wire       [1:0]    _zz_17;
  wire       [1:0]    _zz_18;
  wire       [1:0]    _zz_19;
  wire       [1:0]    _zz_20;
  wire       [1:0]    _zz_21;
  wire       [1:0]    _zz_22;
  wire       [1:0]    _zz_23;
  wire       [1:0]    _zz_24;
  wire       [1:0]    _zz_25;
  wire       [1:0]    _zz_26;
  wire       [1:0]    _zz_27;
  wire       [1:0]    _zz_28;
  wire       [1:0]    _zz_29;
  wire       [1:0]    _zz_30;
  wire       [1:0]    _zz_31;
  wire       [1:0]    _zz_32;
  wire       [1:0]    _zz_33;
  wire       [1:0]    _zz_34;
  wire       [1:0]    _zz_35;
  wire       [1:0]    _zz_36;
  wire       [1:0]    _zz_37;
  wire       [1:0]    _zz_38;
  wire       [1:0]    _zz_39;
  wire       [1:0]    _zz_40;
  wire       [1:0]    _zz_41;
  wire       [1:0]    _zz_42;
  wire       [1:0]    _zz_43;
  wire       [1:0]    _zz_44;
  wire       [1:0]    _zz_45;
  wire       [1:0]    _zz_46;
  wire       [1:0]    _zz_47;
  wire       [1:0]    _zz_48;
  wire       [1:0]    _zz_49;
  wire       [1:0]    _zz_50;
  wire       [1:0]    _zz_51;
  wire       [1:0]    _zz_52;
  wire       [1:0]    _zz_53;
  wire       [1:0]    _zz_54;
  wire       [1:0]    _zz_55;
  wire       [1:0]    _zz_56;
  wire       [1:0]    _zz_57;
  wire       [1:0]    _zz_58;
  wire       [1:0]    _zz_59;
  wire       [1:0]    _zz_60;
  wire       [1:0]    _zz_61;
  wire       [1:0]    _zz_62;
  wire       [1:0]    _zz_63;
  wire       [1:0]    _zz_64;
  wire       [1:0]    _zz_65;
  wire       [1:0]    _zz_66;
  wire       [1:0]    _zz_67;
  wire       [1:0]    _zz_68;
  wire       [1:0]    _zz_69;
  wire       [1:0]    _zz_70;
  wire       [1:0]    _zz_71;
  wire       [1:0]    _zz_72;
  wire       [1:0]    _zz_73;
  wire       [1:0]    _zz_74;
  wire       [1:0]    _zz_75;
  wire       [1:0]    _zz_76;
  wire       [1:0]    _zz_77;
  wire       [1:0]    _zz_78;
  wire       [1:0]    _zz_79;
  wire       [1:0]    _zz_80;
  wire       [1:0]    _zz_81;
  wire       [1:0]    _zz_82;
  wire       [1:0]    _zz_83;
  wire       [1:0]    _zz_84;
  wire       [1:0]    _zz_85;
  wire       [1:0]    _zz_86;
  wire       [1:0]    _zz_87;
  wire       [1:0]    _zz_88;
  wire       [1:0]    _zz_89;
  wire       [1:0]    _zz_90;
  wire       [1:0]    _zz_91;
  wire       [1:0]    _zz_92;
  wire       [1:0]    _zz_93;
  wire       [1:0]    _zz_94;
  wire       [1:0]    _zz_95;
  wire       [1:0]    _zz_96;
  wire       [1:0]    _zz_97;
  wire       [1:0]    _zz_98;
  wire       [1:0]    _zz_99;
  wire       [1:0]    _zz_100;
  wire       [1:0]    _zz_101;
  wire       [1:0]    _zz_102;
  wire       [1:0]    _zz_103;
  reg        [6:0]    idxLatch;
  reg                 staLatch;
  wire                machine_wantExit;
  reg                 machine_wantStart;
  reg        `machine_enumDefinition_1_defaultEncoding_type machine_stateReg;
  reg        `machine_enumDefinition_1_defaultEncoding_type machine_stateNext;
  `ifndef SYNTHESIS
  reg [127:0] machine_stateReg_string;
  reg [127:0] machine_stateNext_string;
  `endif

  (* ram_init_file = "../VerilogHDL/hid.mif" *) reg [7:0] hidKeyTable [0:127];

  assign _zz_115 = _zz_1[0 : 0];
  assign _zz_116 = _zz_1[1 : 1];
  assign _zz_117 = _zz_2[0 : 0];
  assign _zz_118 = _zz_2[1 : 1];
  assign _zz_119 = _zz_3[0 : 0];
  assign _zz_120 = _zz_3[1 : 1];
  assign _zz_121 = _zz_4[0 : 0];
  assign _zz_122 = _zz_4[1 : 1];
  assign _zz_123 = _zz_5[0 : 0];
  assign _zz_124 = _zz_5[1 : 1];
  assign _zz_125 = _zz_6[0 : 0];
  assign _zz_126 = _zz_6[1 : 1];
  assign _zz_127 = _zz_7[0 : 0];
  assign _zz_128 = _zz_7[1 : 1];
  assign _zz_129 = _zz_8[0 : 0];
  assign _zz_130 = _zz_8[1 : 1];
  assign _zz_131 = _zz_9[0 : 0];
  assign _zz_132 = _zz_9[1 : 1];
  assign _zz_133 = _zz_10[0 : 0];
  assign _zz_134 = _zz_10[1 : 1];
  assign _zz_135 = _zz_11[0 : 0];
  assign _zz_136 = _zz_11[1 : 1];
  assign _zz_137 = _zz_12[0 : 0];
  assign _zz_138 = _zz_12[1 : 1];
  assign _zz_139 = _zz_13[0 : 0];
  assign _zz_140 = _zz_13[1 : 1];
  assign _zz_141 = _zz_14[0 : 0];
  assign _zz_142 = _zz_14[1 : 1];
  assign _zz_143 = _zz_15[0 : 0];
  assign _zz_144 = _zz_15[1 : 1];
  assign _zz_145 = _zz_16[0 : 0];
  assign _zz_146 = _zz_16[1 : 1];
  assign _zz_147 = _zz_17[0 : 0];
  assign _zz_148 = _zz_17[1 : 1];
  assign _zz_149 = _zz_18[0 : 0];
  assign _zz_150 = _zz_18[1 : 1];
  assign _zz_151 = _zz_19[0 : 0];
  assign _zz_152 = _zz_19[1 : 1];
  assign _zz_153 = _zz_20[0 : 0];
  assign _zz_154 = _zz_20[1 : 1];
  assign _zz_155 = _zz_21[0 : 0];
  assign _zz_156 = _zz_21[1 : 1];
  assign _zz_157 = _zz_22[0 : 0];
  assign _zz_158 = _zz_22[1 : 1];
  assign _zz_159 = _zz_23[0 : 0];
  assign _zz_160 = _zz_23[1 : 1];
  assign _zz_161 = _zz_24[0 : 0];
  assign _zz_162 = _zz_24[1 : 1];
  assign _zz_163 = _zz_25[0 : 0];
  assign _zz_164 = _zz_25[1 : 1];
  assign _zz_165 = _zz_26[0 : 0];
  assign _zz_166 = _zz_26[1 : 1];
  assign _zz_167 = _zz_27[0 : 0];
  assign _zz_168 = _zz_27[1 : 1];
  assign _zz_169 = _zz_28[0 : 0];
  assign _zz_170 = _zz_28[1 : 1];
  assign _zz_171 = _zz_29[0 : 0];
  assign _zz_172 = _zz_29[1 : 1];
  assign _zz_173 = _zz_30[0 : 0];
  assign _zz_174 = _zz_30[1 : 1];
  assign _zz_175 = _zz_31[0 : 0];
  assign _zz_176 = _zz_31[1 : 1];
  assign _zz_177 = _zz_32[0 : 0];
  assign _zz_178 = _zz_32[1 : 1];
  assign _zz_179 = _zz_33[0 : 0];
  assign _zz_180 = _zz_33[1 : 1];
  assign _zz_181 = _zz_34[0 : 0];
  assign _zz_182 = _zz_34[1 : 1];
  assign _zz_183 = _zz_35[0 : 0];
  assign _zz_184 = _zz_35[1 : 1];
  assign _zz_185 = _zz_36[0 : 0];
  assign _zz_186 = _zz_36[1 : 1];
  assign _zz_187 = _zz_37[0 : 0];
  assign _zz_188 = _zz_37[1 : 1];
  assign _zz_189 = _zz_38[0 : 0];
  assign _zz_190 = _zz_38[1 : 1];
  assign _zz_191 = _zz_39[0 : 0];
  assign _zz_192 = _zz_39[1 : 1];
  assign _zz_193 = _zz_40[0 : 0];
  assign _zz_194 = _zz_40[1 : 1];
  assign _zz_195 = _zz_41[0 : 0];
  assign _zz_196 = _zz_41[1 : 1];
  assign _zz_197 = _zz_42[0 : 0];
  assign _zz_198 = _zz_42[1 : 1];
  assign _zz_199 = _zz_43[0 : 0];
  assign _zz_200 = _zz_43[1 : 1];
  assign _zz_201 = _zz_44[0 : 0];
  assign _zz_202 = _zz_44[1 : 1];
  assign _zz_203 = _zz_45[0 : 0];
  assign _zz_204 = _zz_45[1 : 1];
  assign _zz_205 = _zz_46[0 : 0];
  assign _zz_206 = _zz_46[1 : 1];
  assign _zz_207 = _zz_47[0 : 0];
  assign _zz_208 = _zz_47[1 : 1];
  assign _zz_209 = _zz_48[0 : 0];
  assign _zz_210 = _zz_48[1 : 1];
  assign _zz_211 = _zz_49[0 : 0];
  assign _zz_212 = _zz_49[1 : 1];
  assign _zz_213 = _zz_50[0 : 0];
  assign _zz_214 = _zz_50[1 : 1];
  assign _zz_215 = _zz_51[0 : 0];
  assign _zz_216 = _zz_51[1 : 1];
  assign _zz_217 = _zz_52[0 : 0];
  assign _zz_218 = _zz_52[1 : 1];
  assign _zz_219 = _zz_53[0 : 0];
  assign _zz_220 = _zz_53[1 : 1];
  assign _zz_221 = _zz_54[0 : 0];
  assign _zz_222 = _zz_54[1 : 1];
  assign _zz_223 = _zz_55[0 : 0];
  assign _zz_224 = _zz_55[1 : 1];
  assign _zz_225 = _zz_56[0 : 0];
  assign _zz_226 = _zz_56[1 : 1];
  assign _zz_227 = _zz_57[0 : 0];
  assign _zz_228 = _zz_57[1 : 1];
  assign _zz_229 = _zz_58[0 : 0];
  assign _zz_230 = _zz_58[1 : 1];
  assign _zz_231 = _zz_59[0 : 0];
  assign _zz_232 = _zz_59[1 : 1];
  assign _zz_233 = _zz_60[0 : 0];
  assign _zz_234 = _zz_60[1 : 1];
  assign _zz_235 = _zz_61[0 : 0];
  assign _zz_236 = _zz_61[1 : 1];
  assign _zz_237 = _zz_62[0 : 0];
  assign _zz_238 = _zz_62[1 : 1];
  assign _zz_239 = _zz_63[0 : 0];
  assign _zz_240 = _zz_63[1 : 1];
  assign _zz_241 = _zz_64[0 : 0];
  assign _zz_242 = _zz_64[1 : 1];
  assign _zz_243 = _zz_65[0 : 0];
  assign _zz_244 = _zz_65[1 : 1];
  assign _zz_245 = _zz_66[0 : 0];
  assign _zz_246 = _zz_66[1 : 1];
  assign _zz_247 = _zz_67[0 : 0];
  assign _zz_248 = _zz_67[1 : 1];
  assign _zz_249 = _zz_68[0 : 0];
  assign _zz_250 = _zz_68[1 : 1];
  assign _zz_251 = _zz_69[0 : 0];
  assign _zz_252 = _zz_69[1 : 1];
  assign _zz_253 = _zz_70[0 : 0];
  assign _zz_254 = _zz_70[1 : 1];
  assign _zz_255 = _zz_71[0 : 0];
  assign _zz_256 = _zz_71[1 : 1];
  assign _zz_257 = _zz_72[0 : 0];
  assign _zz_258 = _zz_72[1 : 1];
  assign _zz_259 = _zz_73[0 : 0];
  assign _zz_260 = _zz_73[1 : 1];
  assign _zz_261 = _zz_74[0 : 0];
  assign _zz_262 = _zz_74[1 : 1];
  assign _zz_263 = _zz_75[0 : 0];
  assign _zz_264 = _zz_75[1 : 1];
  assign _zz_265 = _zz_76[0 : 0];
  assign _zz_266 = _zz_76[1 : 1];
  assign _zz_267 = _zz_77[0 : 0];
  assign _zz_268 = _zz_77[1 : 1];
  assign _zz_269 = _zz_78[0 : 0];
  assign _zz_270 = _zz_78[1 : 1];
  assign _zz_271 = _zz_79[0 : 0];
  assign _zz_272 = _zz_79[1 : 1];
  assign _zz_273 = _zz_80[0 : 0];
  assign _zz_274 = _zz_80[1 : 1];
  assign _zz_275 = _zz_81[0 : 0];
  assign _zz_276 = _zz_81[1 : 1];
  assign _zz_277 = _zz_82[0 : 0];
  assign _zz_278 = _zz_82[1 : 1];
  assign _zz_279 = _zz_83[0 : 0];
  assign _zz_280 = _zz_83[1 : 1];
  assign _zz_281 = _zz_84[0 : 0];
  assign _zz_282 = _zz_84[1 : 1];
  assign _zz_283 = _zz_85[0 : 0];
  assign _zz_284 = _zz_85[1 : 1];
  assign _zz_285 = _zz_86[0 : 0];
  assign _zz_286 = _zz_86[1 : 1];
  assign _zz_287 = _zz_87[0 : 0];
  assign _zz_288 = _zz_87[1 : 1];
  assign _zz_289 = _zz_88[0 : 0];
  assign _zz_290 = _zz_88[1 : 1];
  assign _zz_291 = _zz_89[0 : 0];
  assign _zz_292 = _zz_89[1 : 1];
  assign _zz_293 = _zz_90[0 : 0];
  assign _zz_294 = _zz_90[1 : 1];
  assign _zz_295 = _zz_91[0 : 0];
  assign _zz_296 = _zz_91[1 : 1];
  assign _zz_297 = _zz_92[0 : 0];
  assign _zz_298 = _zz_92[1 : 1];
  assign _zz_299 = _zz_93[0 : 0];
  assign _zz_300 = _zz_93[1 : 1];
  assign _zz_301 = _zz_94[0 : 0];
  assign _zz_302 = _zz_94[1 : 1];
  assign _zz_303 = _zz_95[0 : 0];
  assign _zz_304 = _zz_95[1 : 1];
  assign _zz_305 = _zz_96[0 : 0];
  assign _zz_306 = _zz_96[1 : 1];
  assign _zz_307 = _zz_97[0 : 0];
  assign _zz_308 = _zz_97[1 : 1];
  assign _zz_309 = _zz_98[0 : 0];
  assign _zz_310 = _zz_98[1 : 1];
  assign _zz_311 = _zz_99[0 : 0];
  assign _zz_312 = _zz_99[1 : 1];
  assign _zz_313 = _zz_100[0 : 0];
  assign _zz_314 = _zz_100[1 : 1];
  assign _zz_315 = _zz_101[0 : 0];
  assign _zz_316 = _zz_101[1 : 1];
  assign _zz_317 = _zz_102[0 : 0];
  assign _zz_318 = _zz_102[1 : 1];
  assign _zz_319 = _zz_103[0 : 0];
  assign _zz_320 = _zz_103[1 : 1];
  assign _zz_321 = 1'b1;
  always @ (posedge CLK_50) begin
    if(_zz_321) begin
      _zz_114 <= hidKeyTable[idxLatch];
    end
  end

  UartCtrl uartCtrl_1 (
    .io_config_frame_dataLength    (_zz_105[2:0]                     ), //i
    .io_config_frame_stop          (_zz_106                          ), //i
    .io_config_frame_parity        (_zz_107[1:0]                     ), //i
    .io_config_clockDivider        (_zz_108[19:0]                    ), //i
    .io_write_valid                (_zz_109                          ), //i
    .io_write_ready                (uartCtrl_1_io_write_ready        ), //o
    .io_write_payload              (_zz_110[7:0]                     ), //i
    .io_read_valid                 (uartCtrl_1_io_read_valid         ), //o
    .io_read_ready                 (_zz_111                          ), //i
    .io_read_payload               (uartCtrl_1_io_read_payload[7:0]  ), //o
    .io_uart_txd                   (uartCtrl_1_io_uart_txd           ), //o
    .io_uart_rxd                   (_zz_112                          ), //i
    .io_readError                  (uartCtrl_1_io_readError          ), //o
    .io_writeBreak                 (_zz_113                          ), //i
    .io_readBreak                  (uartCtrl_1_io_readBreak          ), //o
    .CLK_50                        (CLK_50                           ), //i
    ._zz_1                         (_zz_104                          )  //i
  );
  `ifndef SYNTHESIS
  always @(*) begin
    case(machine_stateReg)
      `machine_enumDefinition_1_defaultEncoding_machine_BOOT : machine_stateReg_string = "machine_BOOT    ";
      `machine_enumDefinition_1_defaultEncoding_machine_idle : machine_stateReg_string = "machine_idle    ";
      `machine_enumDefinition_1_defaultEncoding_machine_k6 : machine_stateReg_string = "machine_k6      ";
      `machine_enumDefinition_1_defaultEncoding_machine_k5 : machine_stateReg_string = "machine_k5      ";
      `machine_enumDefinition_1_defaultEncoding_machine_k4 : machine_stateReg_string = "machine_k4      ";
      `machine_enumDefinition_1_defaultEncoding_machine_k3 : machine_stateReg_string = "machine_k3      ";
      `machine_enumDefinition_1_defaultEncoding_machine_k2 : machine_stateReg_string = "machine_k2      ";
      `machine_enumDefinition_1_defaultEncoding_machine_k1 : machine_stateReg_string = "machine_k1      ";
      `machine_enumDefinition_1_defaultEncoding_machine_reserved : machine_stateReg_string = "machine_reserved";
      `machine_enumDefinition_1_defaultEncoding_machine_special : machine_stateReg_string = "machine_special ";
      default : machine_stateReg_string = "????????????????";
    endcase
  end
  always @(*) begin
    case(machine_stateNext)
      `machine_enumDefinition_1_defaultEncoding_machine_BOOT : machine_stateNext_string = "machine_BOOT    ";
      `machine_enumDefinition_1_defaultEncoding_machine_idle : machine_stateNext_string = "machine_idle    ";
      `machine_enumDefinition_1_defaultEncoding_machine_k6 : machine_stateNext_string = "machine_k6      ";
      `machine_enumDefinition_1_defaultEncoding_machine_k5 : machine_stateNext_string = "machine_k5      ";
      `machine_enumDefinition_1_defaultEncoding_machine_k4 : machine_stateNext_string = "machine_k4      ";
      `machine_enumDefinition_1_defaultEncoding_machine_k3 : machine_stateNext_string = "machine_k3      ";
      `machine_enumDefinition_1_defaultEncoding_machine_k2 : machine_stateNext_string = "machine_k2      ";
      `machine_enumDefinition_1_defaultEncoding_machine_k1 : machine_stateNext_string = "machine_k1      ";
      `machine_enumDefinition_1_defaultEncoding_machine_reserved : machine_stateNext_string = "machine_reserved";
      `machine_enumDefinition_1_defaultEncoding_machine_special : machine_stateNext_string = "machine_special ";
      default : machine_stateNext_string = "????????????????";
    endcase
  end
  `endif

  assign _zz_1 = keyBits[1 : 0];
  assign keyStatus_0_valid = _zz_115[0];
  assign keyStatus_0_payload = _zz_116[0];
  assign _zz_2 = keyBits[3 : 2];
  assign keyStatus_1_valid = _zz_117[0];
  assign keyStatus_1_payload = _zz_118[0];
  assign _zz_3 = keyBits[5 : 4];
  assign keyStatus_2_valid = _zz_119[0];
  assign keyStatus_2_payload = _zz_120[0];
  assign _zz_4 = keyBits[7 : 6];
  assign keyStatus_3_valid = _zz_121[0];
  assign keyStatus_3_payload = _zz_122[0];
  assign _zz_5 = keyBits[9 : 8];
  assign keyStatus_4_valid = _zz_123[0];
  assign keyStatus_4_payload = _zz_124[0];
  assign _zz_6 = keyBits[11 : 10];
  assign keyStatus_5_valid = _zz_125[0];
  assign keyStatus_5_payload = _zz_126[0];
  assign _zz_7 = keyBits[13 : 12];
  assign keyStatus_6_valid = _zz_127[0];
  assign keyStatus_6_payload = _zz_128[0];
  assign _zz_8 = keyBits[15 : 14];
  assign keyStatus_7_valid = _zz_129[0];
  assign keyStatus_7_payload = _zz_130[0];
  assign _zz_9 = keyBits[17 : 16];
  assign keyStatus_8_valid = _zz_131[0];
  assign keyStatus_8_payload = _zz_132[0];
  assign _zz_10 = keyBits[19 : 18];
  assign keyStatus_9_valid = _zz_133[0];
  assign keyStatus_9_payload = _zz_134[0];
  assign _zz_11 = keyBits[21 : 20];
  assign keyStatus_10_valid = _zz_135[0];
  assign keyStatus_10_payload = _zz_136[0];
  assign _zz_12 = keyBits[23 : 22];
  assign keyStatus_11_valid = _zz_137[0];
  assign keyStatus_11_payload = _zz_138[0];
  assign _zz_13 = keyBits[25 : 24];
  assign keyStatus_12_valid = _zz_139[0];
  assign keyStatus_12_payload = _zz_140[0];
  assign _zz_14 = keyBits[27 : 26];
  assign keyStatus_13_valid = _zz_141[0];
  assign keyStatus_13_payload = _zz_142[0];
  assign _zz_15 = keyBits[29 : 28];
  assign keyStatus_14_valid = _zz_143[0];
  assign keyStatus_14_payload = _zz_144[0];
  assign _zz_16 = keyBits[31 : 30];
  assign keyStatus_15_valid = _zz_145[0];
  assign keyStatus_15_payload = _zz_146[0];
  assign _zz_17 = keyBits[33 : 32];
  assign keyStatus_16_valid = _zz_147[0];
  assign keyStatus_16_payload = _zz_148[0];
  assign _zz_18 = keyBits[35 : 34];
  assign keyStatus_17_valid = _zz_149[0];
  assign keyStatus_17_payload = _zz_150[0];
  assign _zz_19 = keyBits[37 : 36];
  assign keyStatus_18_valid = _zz_151[0];
  assign keyStatus_18_payload = _zz_152[0];
  assign _zz_20 = keyBits[39 : 38];
  assign keyStatus_19_valid = _zz_153[0];
  assign keyStatus_19_payload = _zz_154[0];
  assign _zz_21 = keyBits[41 : 40];
  assign keyStatus_20_valid = _zz_155[0];
  assign keyStatus_20_payload = _zz_156[0];
  assign _zz_22 = keyBits[43 : 42];
  assign keyStatus_21_valid = _zz_157[0];
  assign keyStatus_21_payload = _zz_158[0];
  assign _zz_23 = keyBits[45 : 44];
  assign keyStatus_22_valid = _zz_159[0];
  assign keyStatus_22_payload = _zz_160[0];
  assign _zz_24 = keyBits[47 : 46];
  assign keyStatus_23_valid = _zz_161[0];
  assign keyStatus_23_payload = _zz_162[0];
  assign _zz_25 = keyBits[49 : 48];
  assign keyStatus_24_valid = _zz_163[0];
  assign keyStatus_24_payload = _zz_164[0];
  assign _zz_26 = keyBits[51 : 50];
  assign keyStatus_25_valid = _zz_165[0];
  assign keyStatus_25_payload = _zz_166[0];
  assign _zz_27 = keyBits[53 : 52];
  assign keyStatus_26_valid = _zz_167[0];
  assign keyStatus_26_payload = _zz_168[0];
  assign _zz_28 = keyBits[55 : 54];
  assign keyStatus_27_valid = _zz_169[0];
  assign keyStatus_27_payload = _zz_170[0];
  assign _zz_29 = keyBits[57 : 56];
  assign keyStatus_28_valid = _zz_171[0];
  assign keyStatus_28_payload = _zz_172[0];
  assign _zz_30 = keyBits[59 : 58];
  assign keyStatus_29_valid = _zz_173[0];
  assign keyStatus_29_payload = _zz_174[0];
  assign _zz_31 = keyBits[61 : 60];
  assign keyStatus_30_valid = _zz_175[0];
  assign keyStatus_30_payload = _zz_176[0];
  assign _zz_32 = keyBits[63 : 62];
  assign keyStatus_31_valid = _zz_177[0];
  assign keyStatus_31_payload = _zz_178[0];
  assign _zz_33 = keyBits[65 : 64];
  assign keyStatus_32_valid = _zz_179[0];
  assign keyStatus_32_payload = _zz_180[0];
  assign _zz_34 = keyBits[67 : 66];
  assign keyStatus_33_valid = _zz_181[0];
  assign keyStatus_33_payload = _zz_182[0];
  assign _zz_35 = keyBits[69 : 68];
  assign keyStatus_34_valid = _zz_183[0];
  assign keyStatus_34_payload = _zz_184[0];
  assign _zz_36 = keyBits[71 : 70];
  assign keyStatus_35_valid = _zz_185[0];
  assign keyStatus_35_payload = _zz_186[0];
  assign _zz_37 = keyBits[73 : 72];
  assign keyStatus_36_valid = _zz_187[0];
  assign keyStatus_36_payload = _zz_188[0];
  assign _zz_38 = keyBits[75 : 74];
  assign keyStatus_37_valid = _zz_189[0];
  assign keyStatus_37_payload = _zz_190[0];
  assign _zz_39 = keyBits[77 : 76];
  assign keyStatus_38_valid = _zz_191[0];
  assign keyStatus_38_payload = _zz_192[0];
  assign _zz_40 = keyBits[79 : 78];
  assign keyStatus_39_valid = _zz_193[0];
  assign keyStatus_39_payload = _zz_194[0];
  assign _zz_41 = keyBits[81 : 80];
  assign keyStatus_40_valid = _zz_195[0];
  assign keyStatus_40_payload = _zz_196[0];
  assign _zz_42 = keyBits[83 : 82];
  assign keyStatus_41_valid = _zz_197[0];
  assign keyStatus_41_payload = _zz_198[0];
  assign _zz_43 = keyBits[85 : 84];
  assign keyStatus_42_valid = _zz_199[0];
  assign keyStatus_42_payload = _zz_200[0];
  assign _zz_44 = keyBits[87 : 86];
  assign keyStatus_43_valid = _zz_201[0];
  assign keyStatus_43_payload = _zz_202[0];
  assign _zz_45 = keyBits[89 : 88];
  assign keyStatus_44_valid = _zz_203[0];
  assign keyStatus_44_payload = _zz_204[0];
  assign _zz_46 = keyBits[91 : 90];
  assign keyStatus_45_valid = _zz_205[0];
  assign keyStatus_45_payload = _zz_206[0];
  assign _zz_47 = keyBits[93 : 92];
  assign keyStatus_46_valid = _zz_207[0];
  assign keyStatus_46_payload = _zz_208[0];
  assign _zz_48 = keyBits[95 : 94];
  assign keyStatus_47_valid = _zz_209[0];
  assign keyStatus_47_payload = _zz_210[0];
  assign _zz_49 = keyBits[97 : 96];
  assign keyStatus_48_valid = _zz_211[0];
  assign keyStatus_48_payload = _zz_212[0];
  assign _zz_50 = keyBits[99 : 98];
  assign keyStatus_49_valid = _zz_213[0];
  assign keyStatus_49_payload = _zz_214[0];
  assign _zz_51 = keyBits[101 : 100];
  assign keyStatus_50_valid = _zz_215[0];
  assign keyStatus_50_payload = _zz_216[0];
  assign _zz_52 = keyBits[103 : 102];
  assign keyStatus_51_valid = _zz_217[0];
  assign keyStatus_51_payload = _zz_218[0];
  assign _zz_53 = keyBits[105 : 104];
  assign keyStatus_52_valid = _zz_219[0];
  assign keyStatus_52_payload = _zz_220[0];
  assign _zz_54 = keyBits[107 : 106];
  assign keyStatus_53_valid = _zz_221[0];
  assign keyStatus_53_payload = _zz_222[0];
  assign _zz_55 = keyBits[109 : 108];
  assign keyStatus_54_valid = _zz_223[0];
  assign keyStatus_54_payload = _zz_224[0];
  assign _zz_56 = keyBits[111 : 110];
  assign keyStatus_55_valid = _zz_225[0];
  assign keyStatus_55_payload = _zz_226[0];
  assign _zz_57 = keyBits[113 : 112];
  assign keyStatus_56_valid = _zz_227[0];
  assign keyStatus_56_payload = _zz_228[0];
  assign _zz_58 = keyBits[115 : 114];
  assign keyStatus_57_valid = _zz_229[0];
  assign keyStatus_57_payload = _zz_230[0];
  assign _zz_59 = keyBits[117 : 116];
  assign keyStatus_58_valid = _zz_231[0];
  assign keyStatus_58_payload = _zz_232[0];
  assign _zz_60 = keyBits[119 : 118];
  assign keyStatus_59_valid = _zz_233[0];
  assign keyStatus_59_payload = _zz_234[0];
  assign _zz_61 = keyBits[121 : 120];
  assign keyStatus_60_valid = _zz_235[0];
  assign keyStatus_60_payload = _zz_236[0];
  assign _zz_62 = keyBits[123 : 122];
  assign keyStatus_61_valid = _zz_237[0];
  assign keyStatus_61_payload = _zz_238[0];
  assign _zz_63 = keyBits[125 : 124];
  assign keyStatus_62_valid = _zz_239[0];
  assign keyStatus_62_payload = _zz_240[0];
  assign _zz_64 = keyBits[127 : 126];
  assign keyStatus_63_valid = _zz_241[0];
  assign keyStatus_63_payload = _zz_242[0];
  assign _zz_65 = keyBits[129 : 128];
  assign keyStatus_64_valid = _zz_243[0];
  assign keyStatus_64_payload = _zz_244[0];
  assign _zz_66 = keyBits[131 : 130];
  assign keyStatus_65_valid = _zz_245[0];
  assign keyStatus_65_payload = _zz_246[0];
  assign _zz_67 = keyBits[133 : 132];
  assign keyStatus_66_valid = _zz_247[0];
  assign keyStatus_66_payload = _zz_248[0];
  assign _zz_68 = keyBits[135 : 134];
  assign keyStatus_67_valid = _zz_249[0];
  assign keyStatus_67_payload = _zz_250[0];
  assign _zz_69 = keyBits[137 : 136];
  assign keyStatus_68_valid = _zz_251[0];
  assign keyStatus_68_payload = _zz_252[0];
  assign _zz_70 = keyBits[139 : 138];
  assign keyStatus_69_valid = _zz_253[0];
  assign keyStatus_69_payload = _zz_254[0];
  assign _zz_71 = keyBits[141 : 140];
  assign keyStatus_70_valid = _zz_255[0];
  assign keyStatus_70_payload = _zz_256[0];
  assign _zz_72 = keyBits[143 : 142];
  assign keyStatus_71_valid = _zz_257[0];
  assign keyStatus_71_payload = _zz_258[0];
  assign _zz_73 = keyBits[145 : 144];
  assign keyStatus_72_valid = _zz_259[0];
  assign keyStatus_72_payload = _zz_260[0];
  assign _zz_74 = keyBits[147 : 146];
  assign keyStatus_73_valid = _zz_261[0];
  assign keyStatus_73_payload = _zz_262[0];
  assign _zz_75 = keyBits[149 : 148];
  assign keyStatus_74_valid = _zz_263[0];
  assign keyStatus_74_payload = _zz_264[0];
  assign _zz_76 = keyBits[151 : 150];
  assign keyStatus_75_valid = _zz_265[0];
  assign keyStatus_75_payload = _zz_266[0];
  assign _zz_77 = keyBits[153 : 152];
  assign keyStatus_76_valid = _zz_267[0];
  assign keyStatus_76_payload = _zz_268[0];
  assign _zz_78 = keyBits[155 : 154];
  assign keyStatus_77_valid = _zz_269[0];
  assign keyStatus_77_payload = _zz_270[0];
  assign _zz_79 = keyBits[157 : 156];
  assign keyStatus_78_valid = _zz_271[0];
  assign keyStatus_78_payload = _zz_272[0];
  assign _zz_80 = keyBits[159 : 158];
  assign keyStatus_79_valid = _zz_273[0];
  assign keyStatus_79_payload = _zz_274[0];
  assign _zz_81 = keyBits[161 : 160];
  assign keyStatus_80_valid = _zz_275[0];
  assign keyStatus_80_payload = _zz_276[0];
  assign _zz_82 = keyBits[163 : 162];
  assign keyStatus_81_valid = _zz_277[0];
  assign keyStatus_81_payload = _zz_278[0];
  assign _zz_83 = keyBits[165 : 164];
  assign keyStatus_82_valid = _zz_279[0];
  assign keyStatus_82_payload = _zz_280[0];
  assign _zz_84 = keyBits[167 : 166];
  assign keyStatus_83_valid = _zz_281[0];
  assign keyStatus_83_payload = _zz_282[0];
  assign _zz_85 = keyBits[169 : 168];
  assign keyStatus_84_valid = _zz_283[0];
  assign keyStatus_84_payload = _zz_284[0];
  assign _zz_86 = keyBits[171 : 170];
  assign keyStatus_85_valid = _zz_285[0];
  assign keyStatus_85_payload = _zz_286[0];
  assign _zz_87 = keyBits[173 : 172];
  assign keyStatus_86_valid = _zz_287[0];
  assign keyStatus_86_payload = _zz_288[0];
  assign _zz_88 = keyBits[175 : 174];
  assign keyStatus_87_valid = _zz_289[0];
  assign keyStatus_87_payload = _zz_290[0];
  assign _zz_89 = keyBits[177 : 176];
  assign keyStatus_88_valid = _zz_291[0];
  assign keyStatus_88_payload = _zz_292[0];
  assign _zz_90 = keyBits[179 : 178];
  assign keyStatus_89_valid = _zz_293[0];
  assign keyStatus_89_payload = _zz_294[0];
  assign _zz_91 = keyBits[181 : 180];
  assign keyStatus_90_valid = _zz_295[0];
  assign keyStatus_90_payload = _zz_296[0];
  assign _zz_92 = keyBits[183 : 182];
  assign keyStatus_91_valid = _zz_297[0];
  assign keyStatus_91_payload = _zz_298[0];
  assign _zz_93 = keyBits[185 : 184];
  assign keyStatus_92_valid = _zz_299[0];
  assign keyStatus_92_payload = _zz_300[0];
  assign _zz_94 = keyBits[187 : 186];
  assign keyStatus_93_valid = _zz_301[0];
  assign keyStatus_93_payload = _zz_302[0];
  assign _zz_95 = keyBits[189 : 188];
  assign keyStatus_94_valid = _zz_303[0];
  assign keyStatus_94_payload = _zz_304[0];
  assign _zz_96 = keyBits[191 : 190];
  assign keyStatus_95_valid = _zz_305[0];
  assign keyStatus_95_payload = _zz_306[0];
  assign _zz_97 = keyBits[193 : 192];
  assign keyStatus_96_valid = _zz_307[0];
  assign keyStatus_96_payload = _zz_308[0];
  assign _zz_98 = keyBits[195 : 194];
  assign keyStatus_97_valid = _zz_309[0];
  assign keyStatus_97_payload = _zz_310[0];
  assign _zz_99 = keyBits[197 : 196];
  assign keyStatus_98_valid = _zz_311[0];
  assign keyStatus_98_payload = _zz_312[0];
  assign _zz_100 = keyBits[199 : 198];
  assign keyStatus_99_valid = _zz_313[0];
  assign keyStatus_99_payload = _zz_314[0];
  assign _zz_101 = keyBits[201 : 200];
  assign keyStatus_100_valid = _zz_315[0];
  assign keyStatus_100_payload = _zz_316[0];
  assign _zz_102 = keyBits[203 : 202];
  assign keyStatus_101_valid = _zz_317[0];
  assign keyStatus_101_payload = _zz_318[0];
  assign _zz_103 = keyBits[205 : 204];
  assign keyStatus_102_valid = _zz_319[0];
  assign keyStatus_102_payload = _zz_320[0];
  assign _zz_108 = 20'h0028a;
  assign _zz_105 = 3'b111;
  assign _zz_107 = `UartParityType_defaultEncoding_NONE;
  assign _zz_106 = `UartStopType_defaultEncoding_ONE;
  assign _zz_112 = 1'b1;
  assign _zz_113 = 1'b0;
  always @ (*) begin
    _zz_110 = 8'h0;
    case(machine_stateReg)
      `machine_enumDefinition_1_defaultEncoding_machine_idle : begin
      end
      `machine_enumDefinition_1_defaultEncoding_machine_k6 : begin
      end
      `machine_enumDefinition_1_defaultEncoding_machine_k5 : begin
      end
      `machine_enumDefinition_1_defaultEncoding_machine_k4 : begin
      end
      `machine_enumDefinition_1_defaultEncoding_machine_k3 : begin
      end
      `machine_enumDefinition_1_defaultEncoding_machine_k2 : begin
      end
      `machine_enumDefinition_1_defaultEncoding_machine_k1 : begin
        if(staLatch)begin
          _zz_110 = _zz_114;
        end
      end
      `machine_enumDefinition_1_defaultEncoding_machine_reserved : begin
      end
      `machine_enumDefinition_1_defaultEncoding_machine_special : begin
        _zz_110 = {1'b0,{keyStatus_94_payload,{keyStatus_85_payload,{keyStatus_96_payload,{keyStatus_91_payload,{keyStatus_92_payload,{keyStatus_74_payload,keyStatus_90_payload}}}}}}};
      end
      default : begin
      end
    endcase
  end

  assign TXD = uartCtrl_1_io_uart_txd;
  assign machine_wantExit = 1'b0;
  always @ (*) begin
    machine_wantStart = 1'b0;
    case(machine_stateReg)
      `machine_enumDefinition_1_defaultEncoding_machine_idle : begin
      end
      `machine_enumDefinition_1_defaultEncoding_machine_k6 : begin
      end
      `machine_enumDefinition_1_defaultEncoding_machine_k5 : begin
      end
      `machine_enumDefinition_1_defaultEncoding_machine_k4 : begin
      end
      `machine_enumDefinition_1_defaultEncoding_machine_k3 : begin
      end
      `machine_enumDefinition_1_defaultEncoding_machine_k2 : begin
      end
      `machine_enumDefinition_1_defaultEncoding_machine_k1 : begin
      end
      `machine_enumDefinition_1_defaultEncoding_machine_reserved : begin
      end
      `machine_enumDefinition_1_defaultEncoding_machine_special : begin
      end
      default : begin
        machine_wantStart = 1'b1;
      end
    endcase
  end

  assign _zz_109 = (! (machine_stateReg == `machine_enumDefinition_1_defaultEncoding_machine_idle));
  always @ (*) begin
    machine_stateNext = machine_stateReg;
    case(machine_stateReg)
      `machine_enumDefinition_1_defaultEncoding_machine_idle : begin
        if(scanIdx_valid)begin
          machine_stateNext = `machine_enumDefinition_1_defaultEncoding_machine_special;
        end
      end
      `machine_enumDefinition_1_defaultEncoding_machine_k6 : begin
        if(uartCtrl_1_io_write_ready)begin
          machine_stateNext = `machine_enumDefinition_1_defaultEncoding_machine_idle;
        end
      end
      `machine_enumDefinition_1_defaultEncoding_machine_k5 : begin
        if(uartCtrl_1_io_write_ready)begin
          machine_stateNext = `machine_enumDefinition_1_defaultEncoding_machine_k6;
        end
      end
      `machine_enumDefinition_1_defaultEncoding_machine_k4 : begin
        if(uartCtrl_1_io_write_ready)begin
          machine_stateNext = `machine_enumDefinition_1_defaultEncoding_machine_k5;
        end
      end
      `machine_enumDefinition_1_defaultEncoding_machine_k3 : begin
        if(uartCtrl_1_io_write_ready)begin
          machine_stateNext = `machine_enumDefinition_1_defaultEncoding_machine_k4;
        end
      end
      `machine_enumDefinition_1_defaultEncoding_machine_k2 : begin
        if(uartCtrl_1_io_write_ready)begin
          machine_stateNext = `machine_enumDefinition_1_defaultEncoding_machine_k3;
        end
      end
      `machine_enumDefinition_1_defaultEncoding_machine_k1 : begin
        if(uartCtrl_1_io_write_ready)begin
          machine_stateNext = `machine_enumDefinition_1_defaultEncoding_machine_k2;
        end
      end
      `machine_enumDefinition_1_defaultEncoding_machine_reserved : begin
        if(uartCtrl_1_io_write_ready)begin
          machine_stateNext = `machine_enumDefinition_1_defaultEncoding_machine_k1;
        end
      end
      `machine_enumDefinition_1_defaultEncoding_machine_special : begin
        if(uartCtrl_1_io_write_ready)begin
          machine_stateNext = `machine_enumDefinition_1_defaultEncoding_machine_reserved;
        end
      end
      default : begin
      end
    endcase
    if(machine_wantStart)begin
      machine_stateNext = `machine_enumDefinition_1_defaultEncoding_machine_idle;
    end
  end

  always @ (posedge CLK_50 or posedge _zz_104) begin
    if (_zz_104) begin
      idxLatch <= 7'h0;
      staLatch <= 1'b0;
      machine_stateReg <= `machine_enumDefinition_1_defaultEncoding_machine_BOOT;
    end else begin
      if(scanIdx_valid)begin
        idxLatch <= scanIdx_payload[6 : 0];
      end
      if(scanIdx_valid)begin
        staLatch <= scanIdx_payload[7];
      end
      machine_stateReg <= machine_stateNext;
    end
  end


endmodule

module PS2Device (
   inout              PS2_CLK,
   inout              PS2_DAT,
  output reg          receiveFromHost_valid,
  output     [7:0]    receiveFromHost_payload,
  input               sendToHost_valid,
  output reg          sendToHost_ready,
  input      [7:0]    sendToHost_payload,
  input               _zz_3,
  input               CLK_50
);
  reg                 _zz_4;
  reg        [7:0]    _zz_5;
  wire                bus_1_tx_failed;
  wire                bus_1_tx_ready;
  wire                bus_1_rx_valid;
  wire       [7:0]    bus_1_rx_payload;
  reg        [8:0]    _zz_1;
  wire                _zz_2;
  reg                 _zz_2_regNext;
  reg                 ps2ClkArea_clockQuarter;
  reg        [7:0]    tx_buf;
  wire                machine_wantExit;
  reg                 machine_wantStart;
  reg                 bus_1_tx_ready_regNext;
  wire                machine_sending;
  reg        `machine_enumDefinition_defaultEncoding_type machine_stateReg;
  reg        `machine_enumDefinition_defaultEncoding_type machine_stateNext;
  `ifndef SYNTHESIS
  reg [95:0] machine_stateReg_string;
  reg [95:0] machine_stateNext_string;
  `endif


  ps2_bus #(
    .BYTE_DELAY(7'h50) 
  ) bus_1 (
    .clock_quarter    (ps2ClkArea_clockQuarter  ), //i
    .reset            (_zz_3                    ), //i
    .tx_failed        (bus_1_tx_failed          ), //o
    .tx_valid         (_zz_4                    ), //i
    .tx_ready         (bus_1_tx_ready           ), //o
    .tx_payload       (_zz_5[7:0]               ), //i
    .rx_valid         (bus_1_rx_valid           ), //o
    .rx_payload       (bus_1_rx_payload[7:0]    ), //o
    .PS2_CLK          (PS2_CLK                  ), //~
    .PS2_DAT          (PS2_DAT                  )  //~
  );
  `ifndef SYNTHESIS
  always @(*) begin
    case(machine_stateReg)
      `machine_enumDefinition_defaultEncoding_machine_BOOT : machine_stateReg_string = "machine_BOOT";
      `machine_enumDefinition_defaultEncoding_machine_idle : machine_stateReg_string = "machine_idle";
      `machine_enumDefinition_defaultEncoding_machine_init : machine_stateReg_string = "machine_init";
      `machine_enumDefinition_defaultEncoding_machine_tx : machine_stateReg_string = "machine_tx  ";
      `machine_enumDefinition_defaultEncoding_machine_rx : machine_stateReg_string = "machine_rx  ";
      `machine_enumDefinition_defaultEncoding_machine_ack : machine_stateReg_string = "machine_ack ";
      default : machine_stateReg_string = "????????????";
    endcase
  end
  always @(*) begin
    case(machine_stateNext)
      `machine_enumDefinition_defaultEncoding_machine_BOOT : machine_stateNext_string = "machine_BOOT";
      `machine_enumDefinition_defaultEncoding_machine_idle : machine_stateNext_string = "machine_idle";
      `machine_enumDefinition_defaultEncoding_machine_init : machine_stateNext_string = "machine_init";
      `machine_enumDefinition_defaultEncoding_machine_tx : machine_stateNext_string = "machine_tx  ";
      `machine_enumDefinition_defaultEncoding_machine_rx : machine_stateNext_string = "machine_rx  ";
      `machine_enumDefinition_defaultEncoding_machine_ack : machine_stateNext_string = "machine_ack ";
      default : machine_stateNext_string = "????????????";
    endcase
  end
  `endif

  assign _zz_2 = (_zz_1 == 9'h1f3);
  always @ (*) begin
    _zz_4 = 1'b0;
    case(machine_stateReg)
      `machine_enumDefinition_defaultEncoding_machine_idle : begin
        _zz_4 = 1'b0;
      end
      `machine_enumDefinition_defaultEncoding_machine_init : begin
        _zz_4 = 1'b1;
      end
      `machine_enumDefinition_defaultEncoding_machine_tx : begin
        _zz_4 = 1'b1;
      end
      `machine_enumDefinition_defaultEncoding_machine_rx : begin
        _zz_4 = 1'b0;
      end
      `machine_enumDefinition_defaultEncoding_machine_ack : begin
        _zz_4 = 1'b1;
      end
      default : begin
      end
    endcase
  end

  always @ (*) begin
    _zz_5 = 8'h0;
    case(machine_stateReg)
      `machine_enumDefinition_defaultEncoding_machine_idle : begin
      end
      `machine_enumDefinition_defaultEncoding_machine_init : begin
        _zz_5 = 8'haa;
      end
      `machine_enumDefinition_defaultEncoding_machine_tx : begin
        _zz_5 = tx_buf;
      end
      `machine_enumDefinition_defaultEncoding_machine_rx : begin
      end
      `machine_enumDefinition_defaultEncoding_machine_ack : begin
        _zz_5 = 8'hfa;
      end
      default : begin
      end
    endcase
  end

  always @ (*) begin
    sendToHost_ready = 1'b0;
    case(machine_stateReg)
      `machine_enumDefinition_defaultEncoding_machine_idle : begin
        sendToHost_ready = 1'b1;
      end
      `machine_enumDefinition_defaultEncoding_machine_init : begin
      end
      `machine_enumDefinition_defaultEncoding_machine_tx : begin
      end
      `machine_enumDefinition_defaultEncoding_machine_rx : begin
      end
      `machine_enumDefinition_defaultEncoding_machine_ack : begin
      end
      default : begin
      end
    endcase
  end

  assign receiveFromHost_payload = bus_1_rx_payload;
  always @ (*) begin
    receiveFromHost_valid = 1'b0;
    case(machine_stateReg)
      `machine_enumDefinition_defaultEncoding_machine_idle : begin
      end
      `machine_enumDefinition_defaultEncoding_machine_init : begin
      end
      `machine_enumDefinition_defaultEncoding_machine_tx : begin
      end
      `machine_enumDefinition_defaultEncoding_machine_rx : begin
      end
      `machine_enumDefinition_defaultEncoding_machine_ack : begin
        if(machine_sending)begin
          receiveFromHost_valid = 1'b1;
        end
      end
      default : begin
      end
    endcase
  end

  assign machine_wantExit = 1'b0;
  always @ (*) begin
    machine_wantStart = 1'b0;
    case(machine_stateReg)
      `machine_enumDefinition_defaultEncoding_machine_idle : begin
      end
      `machine_enumDefinition_defaultEncoding_machine_init : begin
      end
      `machine_enumDefinition_defaultEncoding_machine_tx : begin
      end
      `machine_enumDefinition_defaultEncoding_machine_rx : begin
      end
      `machine_enumDefinition_defaultEncoding_machine_ack : begin
      end
      default : begin
        machine_wantStart = 1'b1;
      end
    endcase
  end

  assign machine_sending = ((! bus_1_tx_ready) && bus_1_tx_ready_regNext);
  always @ (*) begin
    machine_stateNext = machine_stateReg;
    case(machine_stateReg)
      `machine_enumDefinition_defaultEncoding_machine_idle : begin
        if(sendToHost_valid)begin
          machine_stateNext = `machine_enumDefinition_defaultEncoding_machine_tx;
        end
      end
      `machine_enumDefinition_defaultEncoding_machine_init : begin
        if(((! bus_1_tx_failed) && machine_sending))begin
          machine_stateNext = `machine_enumDefinition_defaultEncoding_machine_idle;
        end
      end
      `machine_enumDefinition_defaultEncoding_machine_tx : begin
        if(machine_sending)begin
          machine_stateNext = `machine_enumDefinition_defaultEncoding_machine_idle;
        end
      end
      `machine_enumDefinition_defaultEncoding_machine_rx : begin
      end
      `machine_enumDefinition_defaultEncoding_machine_ack : begin
        if(machine_sending)begin
          case(bus_1_rx_payload)
            8'hff : begin
              machine_stateNext = `machine_enumDefinition_defaultEncoding_machine_init;
            end
            8'hf3, 8'hed : begin
              machine_stateNext = `machine_enumDefinition_defaultEncoding_machine_rx;
            end
            default : begin
              machine_stateNext = `machine_enumDefinition_defaultEncoding_machine_idle;
            end
          endcase
        end
      end
      default : begin
      end
    endcase
    if(bus_1_rx_valid)begin
      machine_stateNext = `machine_enumDefinition_defaultEncoding_machine_ack;
    end
    if(machine_wantStart)begin
      machine_stateNext = `machine_enumDefinition_defaultEncoding_machine_init;
    end
  end

  always @ (posedge CLK_50 or posedge _zz_3) begin
    if (_zz_3) begin
      _zz_1 <= 9'h0;
      _zz_2_regNext <= 1'b0;
      machine_stateReg <= `machine_enumDefinition_defaultEncoding_machine_BOOT;
    end else begin
      _zz_1 <= (_zz_1 + 9'h001);
      if(_zz_2)begin
        _zz_1 <= 9'h0;
      end
      _zz_2_regNext <= _zz_2;
      machine_stateReg <= machine_stateNext;
    end
  end

  always @ (posedge CLK_50) begin
    if(_zz_2_regNext) begin
      ps2ClkArea_clockQuarter <= (! ps2ClkArea_clockQuarter);
    end
  end

  always @ (posedge CLK_50) begin
    if(sendToHost_valid)begin
      tx_buf <= sendToHost_payload;
    end
    bus_1_tx_ready_regNext <= bus_1_tx_ready;
  end


endmodule

module KeyMatrix (
  input               enabled,
  input      [20:0]   COL,
  output     [5:0]    ROW,
  output              scanIdx_valid,
  output     [7:0]    scanIdx_payload,
  output     [205:0]  keyBits,
  input               _zz_1,
  input               CLK_50
);
  reg                 _zz_9;
  reg                 _zz_10;
  wire       [5:0]    scanK_ROW;
  wire       [102:0]  scanK_key_down;
  wire                debounce_1_keyStatus_0_valid;
  wire                debounce_1_keyStatus_0_payload;
  wire                debounce_1_keyStatus_1_valid;
  wire                debounce_1_keyStatus_1_payload;
  wire                debounce_1_keyStatus_2_valid;
  wire                debounce_1_keyStatus_2_payload;
  wire                debounce_1_keyStatus_3_valid;
  wire                debounce_1_keyStatus_3_payload;
  wire                debounce_1_keyStatus_4_valid;
  wire                debounce_1_keyStatus_4_payload;
  wire                debounce_1_keyStatus_5_valid;
  wire                debounce_1_keyStatus_5_payload;
  wire                debounce_1_keyStatus_6_valid;
  wire                debounce_1_keyStatus_6_payload;
  wire                debounce_1_keyStatus_7_valid;
  wire                debounce_1_keyStatus_7_payload;
  wire                debounce_1_keyStatus_8_valid;
  wire                debounce_1_keyStatus_8_payload;
  wire                debounce_1_keyStatus_9_valid;
  wire                debounce_1_keyStatus_9_payload;
  wire                debounce_1_keyStatus_10_valid;
  wire                debounce_1_keyStatus_10_payload;
  wire                debounce_1_keyStatus_11_valid;
  wire                debounce_1_keyStatus_11_payload;
  wire                debounce_1_keyStatus_12_valid;
  wire                debounce_1_keyStatus_12_payload;
  wire                debounce_1_keyStatus_13_valid;
  wire                debounce_1_keyStatus_13_payload;
  wire                debounce_1_keyStatus_14_valid;
  wire                debounce_1_keyStatus_14_payload;
  wire                debounce_1_keyStatus_15_valid;
  wire                debounce_1_keyStatus_15_payload;
  wire                debounce_1_keyStatus_16_valid;
  wire                debounce_1_keyStatus_16_payload;
  wire                debounce_1_keyStatus_17_valid;
  wire                debounce_1_keyStatus_17_payload;
  wire                debounce_1_keyStatus_18_valid;
  wire                debounce_1_keyStatus_18_payload;
  wire                debounce_1_keyStatus_19_valid;
  wire                debounce_1_keyStatus_19_payload;
  wire                debounce_1_keyStatus_20_valid;
  wire                debounce_1_keyStatus_20_payload;
  wire                debounce_1_keyStatus_21_valid;
  wire                debounce_1_keyStatus_21_payload;
  wire                debounce_1_keyStatus_22_valid;
  wire                debounce_1_keyStatus_22_payload;
  wire                debounce_1_keyStatus_23_valid;
  wire                debounce_1_keyStatus_23_payload;
  wire                debounce_1_keyStatus_24_valid;
  wire                debounce_1_keyStatus_24_payload;
  wire                debounce_1_keyStatus_25_valid;
  wire                debounce_1_keyStatus_25_payload;
  wire                debounce_1_keyStatus_26_valid;
  wire                debounce_1_keyStatus_26_payload;
  wire                debounce_1_keyStatus_27_valid;
  wire                debounce_1_keyStatus_27_payload;
  wire                debounce_1_keyStatus_28_valid;
  wire                debounce_1_keyStatus_28_payload;
  wire                debounce_1_keyStatus_29_valid;
  wire                debounce_1_keyStatus_29_payload;
  wire                debounce_1_keyStatus_30_valid;
  wire                debounce_1_keyStatus_30_payload;
  wire                debounce_1_keyStatus_31_valid;
  wire                debounce_1_keyStatus_31_payload;
  wire                debounce_1_keyStatus_32_valid;
  wire                debounce_1_keyStatus_32_payload;
  wire                debounce_1_keyStatus_33_valid;
  wire                debounce_1_keyStatus_33_payload;
  wire                debounce_1_keyStatus_34_valid;
  wire                debounce_1_keyStatus_34_payload;
  wire                debounce_1_keyStatus_35_valid;
  wire                debounce_1_keyStatus_35_payload;
  wire                debounce_1_keyStatus_36_valid;
  wire                debounce_1_keyStatus_36_payload;
  wire                debounce_1_keyStatus_37_valid;
  wire                debounce_1_keyStatus_37_payload;
  wire                debounce_1_keyStatus_38_valid;
  wire                debounce_1_keyStatus_38_payload;
  wire                debounce_1_keyStatus_39_valid;
  wire                debounce_1_keyStatus_39_payload;
  wire                debounce_1_keyStatus_40_valid;
  wire                debounce_1_keyStatus_40_payload;
  wire                debounce_1_keyStatus_41_valid;
  wire                debounce_1_keyStatus_41_payload;
  wire                debounce_1_keyStatus_42_valid;
  wire                debounce_1_keyStatus_42_payload;
  wire                debounce_1_keyStatus_43_valid;
  wire                debounce_1_keyStatus_43_payload;
  wire                debounce_1_keyStatus_44_valid;
  wire                debounce_1_keyStatus_44_payload;
  wire                debounce_1_keyStatus_45_valid;
  wire                debounce_1_keyStatus_45_payload;
  wire                debounce_1_keyStatus_46_valid;
  wire                debounce_1_keyStatus_46_payload;
  wire                debounce_1_keyStatus_47_valid;
  wire                debounce_1_keyStatus_47_payload;
  wire                debounce_1_keyStatus_48_valid;
  wire                debounce_1_keyStatus_48_payload;
  wire                debounce_1_keyStatus_49_valid;
  wire                debounce_1_keyStatus_49_payload;
  wire                debounce_1_keyStatus_50_valid;
  wire                debounce_1_keyStatus_50_payload;
  wire                debounce_1_keyStatus_51_valid;
  wire                debounce_1_keyStatus_51_payload;
  wire                debounce_1_keyStatus_52_valid;
  wire                debounce_1_keyStatus_52_payload;
  wire                debounce_1_keyStatus_53_valid;
  wire                debounce_1_keyStatus_53_payload;
  wire                debounce_1_keyStatus_54_valid;
  wire                debounce_1_keyStatus_54_payload;
  wire                debounce_1_keyStatus_55_valid;
  wire                debounce_1_keyStatus_55_payload;
  wire                debounce_1_keyStatus_56_valid;
  wire                debounce_1_keyStatus_56_payload;
  wire                debounce_1_keyStatus_57_valid;
  wire                debounce_1_keyStatus_57_payload;
  wire                debounce_1_keyStatus_58_valid;
  wire                debounce_1_keyStatus_58_payload;
  wire                debounce_1_keyStatus_59_valid;
  wire                debounce_1_keyStatus_59_payload;
  wire                debounce_1_keyStatus_60_valid;
  wire                debounce_1_keyStatus_60_payload;
  wire                debounce_1_keyStatus_61_valid;
  wire                debounce_1_keyStatus_61_payload;
  wire                debounce_1_keyStatus_62_valid;
  wire                debounce_1_keyStatus_62_payload;
  wire                debounce_1_keyStatus_63_valid;
  wire                debounce_1_keyStatus_63_payload;
  wire                debounce_1_keyStatus_64_valid;
  wire                debounce_1_keyStatus_64_payload;
  wire                debounce_1_keyStatus_65_valid;
  wire                debounce_1_keyStatus_65_payload;
  wire                debounce_1_keyStatus_66_valid;
  wire                debounce_1_keyStatus_66_payload;
  wire                debounce_1_keyStatus_67_valid;
  wire                debounce_1_keyStatus_67_payload;
  wire                debounce_1_keyStatus_68_valid;
  wire                debounce_1_keyStatus_68_payload;
  wire                debounce_1_keyStatus_69_valid;
  wire                debounce_1_keyStatus_69_payload;
  wire                debounce_1_keyStatus_70_valid;
  wire                debounce_1_keyStatus_70_payload;
  wire                debounce_1_keyStatus_71_valid;
  wire                debounce_1_keyStatus_71_payload;
  wire                debounce_1_keyStatus_72_valid;
  wire                debounce_1_keyStatus_72_payload;
  wire                debounce_1_keyStatus_73_valid;
  wire                debounce_1_keyStatus_73_payload;
  wire                debounce_1_keyStatus_74_valid;
  wire                debounce_1_keyStatus_74_payload;
  wire                debounce_1_keyStatus_75_valid;
  wire                debounce_1_keyStatus_75_payload;
  wire                debounce_1_keyStatus_76_valid;
  wire                debounce_1_keyStatus_76_payload;
  wire                debounce_1_keyStatus_77_valid;
  wire                debounce_1_keyStatus_77_payload;
  wire                debounce_1_keyStatus_78_valid;
  wire                debounce_1_keyStatus_78_payload;
  wire                debounce_1_keyStatus_79_valid;
  wire                debounce_1_keyStatus_79_payload;
  wire                debounce_1_keyStatus_80_valid;
  wire                debounce_1_keyStatus_80_payload;
  wire                debounce_1_keyStatus_81_valid;
  wire                debounce_1_keyStatus_81_payload;
  wire                debounce_1_keyStatus_82_valid;
  wire                debounce_1_keyStatus_82_payload;
  wire                debounce_1_keyStatus_83_valid;
  wire                debounce_1_keyStatus_83_payload;
  wire                debounce_1_keyStatus_84_valid;
  wire                debounce_1_keyStatus_84_payload;
  wire                debounce_1_keyStatus_85_valid;
  wire                debounce_1_keyStatus_85_payload;
  wire                debounce_1_keyStatus_86_valid;
  wire                debounce_1_keyStatus_86_payload;
  wire                debounce_1_keyStatus_87_valid;
  wire                debounce_1_keyStatus_87_payload;
  wire                debounce_1_keyStatus_88_valid;
  wire                debounce_1_keyStatus_88_payload;
  wire                debounce_1_keyStatus_89_valid;
  wire                debounce_1_keyStatus_89_payload;
  wire                debounce_1_keyStatus_90_valid;
  wire                debounce_1_keyStatus_90_payload;
  wire                debounce_1_keyStatus_91_valid;
  wire                debounce_1_keyStatus_91_payload;
  wire                debounce_1_keyStatus_92_valid;
  wire                debounce_1_keyStatus_92_payload;
  wire                debounce_1_keyStatus_93_valid;
  wire                debounce_1_keyStatus_93_payload;
  wire                debounce_1_keyStatus_94_valid;
  wire                debounce_1_keyStatus_94_payload;
  wire                debounce_1_keyStatus_95_valid;
  wire                debounce_1_keyStatus_95_payload;
  wire                debounce_1_keyStatus_96_valid;
  wire                debounce_1_keyStatus_96_payload;
  wire                debounce_1_keyStatus_97_valid;
  wire                debounce_1_keyStatus_97_payload;
  wire                debounce_1_keyStatus_98_valid;
  wire                debounce_1_keyStatus_98_payload;
  wire                debounce_1_keyStatus_99_valid;
  wire                debounce_1_keyStatus_99_payload;
  wire                debounce_1_keyStatus_100_valid;
  wire                debounce_1_keyStatus_100_payload;
  wire                debounce_1_keyStatus_101_valid;
  wire                debounce_1_keyStatus_101_payload;
  wire                debounce_1_keyStatus_102_valid;
  wire                debounce_1_keyStatus_102_payload;
  wire       [0:0]    _zz_11;
  wire       [10:0]   _zz_12;
  wire       [0:0]    _zz_13;
  wire       [6:0]    _zz_14;
  wire       [0:0]    _zz_15;
  wire       [0:0]    _zz_16;
  wire       [1:0]    _zz_17;
  wire       [191:0]  _zz_18;
  wire       [0:0]    _zz_19;
  wire       [0:0]    _zz_20;
  wire       [1:0]    _zz_21;
  wire       [179:0]  _zz_22;
  wire       [0:0]    _zz_23;
  wire       [0:0]    _zz_24;
  wire       [1:0]    _zz_25;
  wire       [167:0]  _zz_26;
  wire       [0:0]    _zz_27;
  wire       [0:0]    _zz_28;
  wire       [1:0]    _zz_29;
  wire       [155:0]  _zz_30;
  wire       [0:0]    _zz_31;
  wire       [0:0]    _zz_32;
  wire       [1:0]    _zz_33;
  wire       [143:0]  _zz_34;
  wire       [0:0]    _zz_35;
  wire       [0:0]    _zz_36;
  wire       [1:0]    _zz_37;
  wire       [131:0]  _zz_38;
  wire       [0:0]    _zz_39;
  wire       [0:0]    _zz_40;
  wire       [1:0]    _zz_41;
  wire       [119:0]  _zz_42;
  wire       [0:0]    _zz_43;
  wire       [0:0]    _zz_44;
  wire       [1:0]    _zz_45;
  wire       [107:0]  _zz_46;
  wire       [0:0]    _zz_47;
  wire       [0:0]    _zz_48;
  wire       [1:0]    _zz_49;
  wire       [95:0]   _zz_50;
  wire       [0:0]    _zz_51;
  wire       [0:0]    _zz_52;
  wire       [1:0]    _zz_53;
  wire       [83:0]   _zz_54;
  wire       [0:0]    _zz_55;
  wire       [0:0]    _zz_56;
  wire       [1:0]    _zz_57;
  wire       [71:0]   _zz_58;
  wire       [0:0]    _zz_59;
  wire       [0:0]    _zz_60;
  wire       [1:0]    _zz_61;
  wire       [59:0]   _zz_62;
  wire       [0:0]    _zz_63;
  wire       [0:0]    _zz_64;
  wire       [1:0]    _zz_65;
  wire       [47:0]   _zz_66;
  wire       [0:0]    _zz_67;
  wire       [0:0]    _zz_68;
  wire       [1:0]    _zz_69;
  wire       [35:0]   _zz_70;
  wire       [0:0]    _zz_71;
  wire       [0:0]    _zz_72;
  wire       [1:0]    _zz_73;
  wire       [23:0]   _zz_74;
  wire       [0:0]    _zz_75;
  wire       [0:0]    _zz_76;
  wire       [1:0]    _zz_77;
  wire       [11:0]   _zz_78;
  wire       [0:0]    _zz_79;
  wire       [0:0]    _zz_80;
  wire       [0:0]    _zz_81;
  wire       [0:0]    _zz_82;
  wire                keyStatus_0_valid;
  wire                keyStatus_0_payload;
  wire                keyStatus_1_valid;
  wire                keyStatus_1_payload;
  wire                keyStatus_2_valid;
  wire                keyStatus_2_payload;
  wire                keyStatus_3_valid;
  wire                keyStatus_3_payload;
  wire                keyStatus_4_valid;
  wire                keyStatus_4_payload;
  wire                keyStatus_5_valid;
  wire                keyStatus_5_payload;
  wire                keyStatus_6_valid;
  wire                keyStatus_6_payload;
  wire                keyStatus_7_valid;
  wire                keyStatus_7_payload;
  wire                keyStatus_8_valid;
  wire                keyStatus_8_payload;
  wire                keyStatus_9_valid;
  wire                keyStatus_9_payload;
  wire                keyStatus_10_valid;
  wire                keyStatus_10_payload;
  wire                keyStatus_11_valid;
  wire                keyStatus_11_payload;
  wire                keyStatus_12_valid;
  wire                keyStatus_12_payload;
  wire                keyStatus_13_valid;
  wire                keyStatus_13_payload;
  wire                keyStatus_14_valid;
  wire                keyStatus_14_payload;
  wire                keyStatus_15_valid;
  wire                keyStatus_15_payload;
  wire                keyStatus_16_valid;
  wire                keyStatus_16_payload;
  wire                keyStatus_17_valid;
  wire                keyStatus_17_payload;
  wire                keyStatus_18_valid;
  wire                keyStatus_18_payload;
  wire                keyStatus_19_valid;
  wire                keyStatus_19_payload;
  wire                keyStatus_20_valid;
  wire                keyStatus_20_payload;
  wire                keyStatus_21_valid;
  wire                keyStatus_21_payload;
  wire                keyStatus_22_valid;
  wire                keyStatus_22_payload;
  wire                keyStatus_23_valid;
  wire                keyStatus_23_payload;
  wire                keyStatus_24_valid;
  wire                keyStatus_24_payload;
  wire                keyStatus_25_valid;
  wire                keyStatus_25_payload;
  wire                keyStatus_26_valid;
  wire                keyStatus_26_payload;
  wire                keyStatus_27_valid;
  wire                keyStatus_27_payload;
  wire                keyStatus_28_valid;
  wire                keyStatus_28_payload;
  wire                keyStatus_29_valid;
  wire                keyStatus_29_payload;
  wire                keyStatus_30_valid;
  wire                keyStatus_30_payload;
  wire                keyStatus_31_valid;
  wire                keyStatus_31_payload;
  wire                keyStatus_32_valid;
  wire                keyStatus_32_payload;
  wire                keyStatus_33_valid;
  wire                keyStatus_33_payload;
  wire                keyStatus_34_valid;
  wire                keyStatus_34_payload;
  wire                keyStatus_35_valid;
  wire                keyStatus_35_payload;
  wire                keyStatus_36_valid;
  wire                keyStatus_36_payload;
  wire                keyStatus_37_valid;
  wire                keyStatus_37_payload;
  wire                keyStatus_38_valid;
  wire                keyStatus_38_payload;
  wire                keyStatus_39_valid;
  wire                keyStatus_39_payload;
  wire                keyStatus_40_valid;
  wire                keyStatus_40_payload;
  wire                keyStatus_41_valid;
  wire                keyStatus_41_payload;
  wire                keyStatus_42_valid;
  wire                keyStatus_42_payload;
  wire                keyStatus_43_valid;
  wire                keyStatus_43_payload;
  wire                keyStatus_44_valid;
  wire                keyStatus_44_payload;
  wire                keyStatus_45_valid;
  wire                keyStatus_45_payload;
  wire                keyStatus_46_valid;
  wire                keyStatus_46_payload;
  wire                keyStatus_47_valid;
  wire                keyStatus_47_payload;
  wire                keyStatus_48_valid;
  wire                keyStatus_48_payload;
  wire                keyStatus_49_valid;
  wire                keyStatus_49_payload;
  wire                keyStatus_50_valid;
  wire                keyStatus_50_payload;
  wire                keyStatus_51_valid;
  wire                keyStatus_51_payload;
  wire                keyStatus_52_valid;
  wire                keyStatus_52_payload;
  wire                keyStatus_53_valid;
  wire                keyStatus_53_payload;
  wire                keyStatus_54_valid;
  wire                keyStatus_54_payload;
  wire                keyStatus_55_valid;
  wire                keyStatus_55_payload;
  wire                keyStatus_56_valid;
  wire                keyStatus_56_payload;
  wire                keyStatus_57_valid;
  wire                keyStatus_57_payload;
  wire                keyStatus_58_valid;
  wire                keyStatus_58_payload;
  wire                keyStatus_59_valid;
  wire                keyStatus_59_payload;
  wire                keyStatus_60_valid;
  wire                keyStatus_60_payload;
  wire                keyStatus_61_valid;
  wire                keyStatus_61_payload;
  wire                keyStatus_62_valid;
  wire                keyStatus_62_payload;
  wire                keyStatus_63_valid;
  wire                keyStatus_63_payload;
  wire                keyStatus_64_valid;
  wire                keyStatus_64_payload;
  wire                keyStatus_65_valid;
  wire                keyStatus_65_payload;
  wire                keyStatus_66_valid;
  wire                keyStatus_66_payload;
  wire                keyStatus_67_valid;
  wire                keyStatus_67_payload;
  wire                keyStatus_68_valid;
  wire                keyStatus_68_payload;
  wire                keyStatus_69_valid;
  wire                keyStatus_69_payload;
  wire                keyStatus_70_valid;
  wire                keyStatus_70_payload;
  wire                keyStatus_71_valid;
  wire                keyStatus_71_payload;
  wire                keyStatus_72_valid;
  wire                keyStatus_72_payload;
  wire                keyStatus_73_valid;
  wire                keyStatus_73_payload;
  wire                keyStatus_74_valid;
  wire                keyStatus_74_payload;
  wire                keyStatus_75_valid;
  wire                keyStatus_75_payload;
  wire                keyStatus_76_valid;
  wire                keyStatus_76_payload;
  wire                keyStatus_77_valid;
  wire                keyStatus_77_payload;
  wire                keyStatus_78_valid;
  wire                keyStatus_78_payload;
  wire                keyStatus_79_valid;
  wire                keyStatus_79_payload;
  wire                keyStatus_80_valid;
  wire                keyStatus_80_payload;
  wire                keyStatus_81_valid;
  wire                keyStatus_81_payload;
  wire                keyStatus_82_valid;
  wire                keyStatus_82_payload;
  wire                keyStatus_83_valid;
  wire                keyStatus_83_payload;
  wire                keyStatus_84_valid;
  wire                keyStatus_84_payload;
  wire                keyStatus_85_valid;
  wire                keyStatus_85_payload;
  wire                keyStatus_86_valid;
  wire                keyStatus_86_payload;
  wire                keyStatus_87_valid;
  wire                keyStatus_87_payload;
  wire                keyStatus_88_valid;
  wire                keyStatus_88_payload;
  wire                keyStatus_89_valid;
  wire                keyStatus_89_payload;
  wire                keyStatus_90_valid;
  wire                keyStatus_90_payload;
  wire                keyStatus_91_valid;
  wire                keyStatus_91_payload;
  wire                keyStatus_92_valid;
  wire                keyStatus_92_payload;
  wire                keyStatus_93_valid;
  wire                keyStatus_93_payload;
  wire                keyStatus_94_valid;
  wire                keyStatus_94_payload;
  wire                keyStatus_95_valid;
  wire                keyStatus_95_payload;
  wire                keyStatus_96_valid;
  wire                keyStatus_96_payload;
  wire                keyStatus_97_valid;
  wire                keyStatus_97_payload;
  wire                keyStatus_98_valid;
  wire                keyStatus_98_payload;
  wire                keyStatus_99_valid;
  wire                keyStatus_99_payload;
  wire                keyStatus_100_valid;
  wire                keyStatus_100_payload;
  wire                keyStatus_101_valid;
  wire                keyStatus_101_payload;
  wire                keyStatus_102_valid;
  wire                keyStatus_102_payload;
  reg                 clkScan_state;
  reg                 clkScan_stateRise;
  wire                clkScan_counter_willIncrement;
  reg                 clkScan_counter_willClear;
  reg        [10:0]   clkScan_counter_valueNext;
  reg        [10:0]   clkScan_counter_value;
  wire                clkScan_counter_willOverflowIfInc;
  wire                clkScan_counter_willOverflow;
  reg        [6:0]    _zz_2;
  wire                _zz_3;
  reg                 _zz_3_regNext;
  wire                _zz_4;
  reg        [6:0]    _zz_5;
  reg        [6:0]    _zz_6;
  wire                _zz_7;
  wire                _zz_8;

  assign _zz_11 = clkScan_counter_willIncrement;
  assign _zz_12 = {10'd0, _zz_11};
  assign _zz_13 = _zz_4;
  assign _zz_14 = {6'd0, _zz_13};
  assign _zz_15 = keyStatus_97_payload;
  assign _zz_16 = keyStatus_97_valid;
  assign _zz_17 = {keyStatus_96_payload,keyStatus_96_valid};
  assign _zz_18 = {{keyStatus_95_payload,keyStatus_95_valid},{{keyStatus_94_payload,keyStatus_94_valid},{{keyStatus_93_payload,keyStatus_93_valid},{{keyStatus_92_payload,keyStatus_92_valid},{{_zz_19,_zz_20},{_zz_21,_zz_22}}}}}};
  assign _zz_19 = keyStatus_91_payload;
  assign _zz_20 = keyStatus_91_valid;
  assign _zz_21 = {keyStatus_90_payload,keyStatus_90_valid};
  assign _zz_22 = {{keyStatus_89_payload,keyStatus_89_valid},{{keyStatus_88_payload,keyStatus_88_valid},{{keyStatus_87_payload,keyStatus_87_valid},{{keyStatus_86_payload,keyStatus_86_valid},{{_zz_23,_zz_24},{_zz_25,_zz_26}}}}}};
  assign _zz_23 = keyStatus_85_payload;
  assign _zz_24 = keyStatus_85_valid;
  assign _zz_25 = {keyStatus_84_payload,keyStatus_84_valid};
  assign _zz_26 = {{keyStatus_83_payload,keyStatus_83_valid},{{keyStatus_82_payload,keyStatus_82_valid},{{keyStatus_81_payload,keyStatus_81_valid},{{keyStatus_80_payload,keyStatus_80_valid},{{_zz_27,_zz_28},{_zz_29,_zz_30}}}}}};
  assign _zz_27 = keyStatus_79_payload;
  assign _zz_28 = keyStatus_79_valid;
  assign _zz_29 = {keyStatus_78_payload,keyStatus_78_valid};
  assign _zz_30 = {{keyStatus_77_payload,keyStatus_77_valid},{{keyStatus_76_payload,keyStatus_76_valid},{{keyStatus_75_payload,keyStatus_75_valid},{{keyStatus_74_payload,keyStatus_74_valid},{{_zz_31,_zz_32},{_zz_33,_zz_34}}}}}};
  assign _zz_31 = keyStatus_73_payload;
  assign _zz_32 = keyStatus_73_valid;
  assign _zz_33 = {keyStatus_72_payload,keyStatus_72_valid};
  assign _zz_34 = {{keyStatus_71_payload,keyStatus_71_valid},{{keyStatus_70_payload,keyStatus_70_valid},{{keyStatus_69_payload,keyStatus_69_valid},{{keyStatus_68_payload,keyStatus_68_valid},{{_zz_35,_zz_36},{_zz_37,_zz_38}}}}}};
  assign _zz_35 = keyStatus_67_payload;
  assign _zz_36 = keyStatus_67_valid;
  assign _zz_37 = {keyStatus_66_payload,keyStatus_66_valid};
  assign _zz_38 = {{keyStatus_65_payload,keyStatus_65_valid},{{keyStatus_64_payload,keyStatus_64_valid},{{keyStatus_63_payload,keyStatus_63_valid},{{keyStatus_62_payload,keyStatus_62_valid},{{_zz_39,_zz_40},{_zz_41,_zz_42}}}}}};
  assign _zz_39 = keyStatus_61_payload;
  assign _zz_40 = keyStatus_61_valid;
  assign _zz_41 = {keyStatus_60_payload,keyStatus_60_valid};
  assign _zz_42 = {{keyStatus_59_payload,keyStatus_59_valid},{{keyStatus_58_payload,keyStatus_58_valid},{{keyStatus_57_payload,keyStatus_57_valid},{{keyStatus_56_payload,keyStatus_56_valid},{{_zz_43,_zz_44},{_zz_45,_zz_46}}}}}};
  assign _zz_43 = keyStatus_55_payload;
  assign _zz_44 = keyStatus_55_valid;
  assign _zz_45 = {keyStatus_54_payload,keyStatus_54_valid};
  assign _zz_46 = {{keyStatus_53_payload,keyStatus_53_valid},{{keyStatus_52_payload,keyStatus_52_valid},{{keyStatus_51_payload,keyStatus_51_valid},{{keyStatus_50_payload,keyStatus_50_valid},{{_zz_47,_zz_48},{_zz_49,_zz_50}}}}}};
  assign _zz_47 = keyStatus_49_payload;
  assign _zz_48 = keyStatus_49_valid;
  assign _zz_49 = {keyStatus_48_payload,keyStatus_48_valid};
  assign _zz_50 = {{keyStatus_47_payload,keyStatus_47_valid},{{keyStatus_46_payload,keyStatus_46_valid},{{keyStatus_45_payload,keyStatus_45_valid},{{keyStatus_44_payload,keyStatus_44_valid},{{_zz_51,_zz_52},{_zz_53,_zz_54}}}}}};
  assign _zz_51 = keyStatus_43_payload;
  assign _zz_52 = keyStatus_43_valid;
  assign _zz_53 = {keyStatus_42_payload,keyStatus_42_valid};
  assign _zz_54 = {{keyStatus_41_payload,keyStatus_41_valid},{{keyStatus_40_payload,keyStatus_40_valid},{{keyStatus_39_payload,keyStatus_39_valid},{{keyStatus_38_payload,keyStatus_38_valid},{{_zz_55,_zz_56},{_zz_57,_zz_58}}}}}};
  assign _zz_55 = keyStatus_37_payload;
  assign _zz_56 = keyStatus_37_valid;
  assign _zz_57 = {keyStatus_36_payload,keyStatus_36_valid};
  assign _zz_58 = {{keyStatus_35_payload,keyStatus_35_valid},{{keyStatus_34_payload,keyStatus_34_valid},{{keyStatus_33_payload,keyStatus_33_valid},{{keyStatus_32_payload,keyStatus_32_valid},{{_zz_59,_zz_60},{_zz_61,_zz_62}}}}}};
  assign _zz_59 = keyStatus_31_payload;
  assign _zz_60 = keyStatus_31_valid;
  assign _zz_61 = {keyStatus_30_payload,keyStatus_30_valid};
  assign _zz_62 = {{keyStatus_29_payload,keyStatus_29_valid},{{keyStatus_28_payload,keyStatus_28_valid},{{keyStatus_27_payload,keyStatus_27_valid},{{keyStatus_26_payload,keyStatus_26_valid},{{_zz_63,_zz_64},{_zz_65,_zz_66}}}}}};
  assign _zz_63 = keyStatus_25_payload;
  assign _zz_64 = keyStatus_25_valid;
  assign _zz_65 = {keyStatus_24_payload,keyStatus_24_valid};
  assign _zz_66 = {{keyStatus_23_payload,keyStatus_23_valid},{{keyStatus_22_payload,keyStatus_22_valid},{{keyStatus_21_payload,keyStatus_21_valid},{{keyStatus_20_payload,keyStatus_20_valid},{{_zz_67,_zz_68},{_zz_69,_zz_70}}}}}};
  assign _zz_67 = keyStatus_19_payload;
  assign _zz_68 = keyStatus_19_valid;
  assign _zz_69 = {keyStatus_18_payload,keyStatus_18_valid};
  assign _zz_70 = {{keyStatus_17_payload,keyStatus_17_valid},{{keyStatus_16_payload,keyStatus_16_valid},{{keyStatus_15_payload,keyStatus_15_valid},{{keyStatus_14_payload,keyStatus_14_valid},{{_zz_71,_zz_72},{_zz_73,_zz_74}}}}}};
  assign _zz_71 = keyStatus_13_payload;
  assign _zz_72 = keyStatus_13_valid;
  assign _zz_73 = {keyStatus_12_payload,keyStatus_12_valid};
  assign _zz_74 = {{keyStatus_11_payload,keyStatus_11_valid},{{keyStatus_10_payload,keyStatus_10_valid},{{keyStatus_9_payload,keyStatus_9_valid},{{keyStatus_8_payload,keyStatus_8_valid},{{_zz_75,_zz_76},{_zz_77,_zz_78}}}}}};
  assign _zz_75 = keyStatus_7_payload;
  assign _zz_76 = keyStatus_7_valid;
  assign _zz_77 = {keyStatus_6_payload,keyStatus_6_valid};
  assign _zz_78 = {{keyStatus_5_payload,keyStatus_5_valid},{{keyStatus_4_payload,keyStatus_4_valid},{{keyStatus_3_payload,keyStatus_3_valid},{{keyStatus_2_payload,keyStatus_2_valid},{{_zz_79,_zz_80},{_zz_81,_zz_82}}}}}};
  assign _zz_79 = keyStatus_1_payload;
  assign _zz_80 = keyStatus_1_valid;
  assign _zz_81 = keyStatus_0_payload;
  assign _zz_82 = keyStatus_0_valid;
  scan_key scanK (
    .clock       (clkScan_state          ), //i
    .reset       (_zz_1                  ), //i
    .enabled     (enabled                ), //i
    .COL         (COL[20:0]              ), //i
    .ROW         (scanK_ROW[5:0]         ), //o
    .key_down    (scanK_key_down[102:0]  )  //o
  );
  Debounce debounce_1 (
    .key_down                 (scanK_key_down[102:0]             ), //i
    .keyStatus_0_valid        (debounce_1_keyStatus_0_valid      ), //o
    .keyStatus_0_payload      (debounce_1_keyStatus_0_payload    ), //o
    .keyStatus_1_valid        (debounce_1_keyStatus_1_valid      ), //o
    .keyStatus_1_payload      (debounce_1_keyStatus_1_payload    ), //o
    .keyStatus_2_valid        (debounce_1_keyStatus_2_valid      ), //o
    .keyStatus_2_payload      (debounce_1_keyStatus_2_payload    ), //o
    .keyStatus_3_valid        (debounce_1_keyStatus_3_valid      ), //o
    .keyStatus_3_payload      (debounce_1_keyStatus_3_payload    ), //o
    .keyStatus_4_valid        (debounce_1_keyStatus_4_valid      ), //o
    .keyStatus_4_payload      (debounce_1_keyStatus_4_payload    ), //o
    .keyStatus_5_valid        (debounce_1_keyStatus_5_valid      ), //o
    .keyStatus_5_payload      (debounce_1_keyStatus_5_payload    ), //o
    .keyStatus_6_valid        (debounce_1_keyStatus_6_valid      ), //o
    .keyStatus_6_payload      (debounce_1_keyStatus_6_payload    ), //o
    .keyStatus_7_valid        (debounce_1_keyStatus_7_valid      ), //o
    .keyStatus_7_payload      (debounce_1_keyStatus_7_payload    ), //o
    .keyStatus_8_valid        (debounce_1_keyStatus_8_valid      ), //o
    .keyStatus_8_payload      (debounce_1_keyStatus_8_payload    ), //o
    .keyStatus_9_valid        (debounce_1_keyStatus_9_valid      ), //o
    .keyStatus_9_payload      (debounce_1_keyStatus_9_payload    ), //o
    .keyStatus_10_valid       (debounce_1_keyStatus_10_valid     ), //o
    .keyStatus_10_payload     (debounce_1_keyStatus_10_payload   ), //o
    .keyStatus_11_valid       (debounce_1_keyStatus_11_valid     ), //o
    .keyStatus_11_payload     (debounce_1_keyStatus_11_payload   ), //o
    .keyStatus_12_valid       (debounce_1_keyStatus_12_valid     ), //o
    .keyStatus_12_payload     (debounce_1_keyStatus_12_payload   ), //o
    .keyStatus_13_valid       (debounce_1_keyStatus_13_valid     ), //o
    .keyStatus_13_payload     (debounce_1_keyStatus_13_payload   ), //o
    .keyStatus_14_valid       (debounce_1_keyStatus_14_valid     ), //o
    .keyStatus_14_payload     (debounce_1_keyStatus_14_payload   ), //o
    .keyStatus_15_valid       (debounce_1_keyStatus_15_valid     ), //o
    .keyStatus_15_payload     (debounce_1_keyStatus_15_payload   ), //o
    .keyStatus_16_valid       (debounce_1_keyStatus_16_valid     ), //o
    .keyStatus_16_payload     (debounce_1_keyStatus_16_payload   ), //o
    .keyStatus_17_valid       (debounce_1_keyStatus_17_valid     ), //o
    .keyStatus_17_payload     (debounce_1_keyStatus_17_payload   ), //o
    .keyStatus_18_valid       (debounce_1_keyStatus_18_valid     ), //o
    .keyStatus_18_payload     (debounce_1_keyStatus_18_payload   ), //o
    .keyStatus_19_valid       (debounce_1_keyStatus_19_valid     ), //o
    .keyStatus_19_payload     (debounce_1_keyStatus_19_payload   ), //o
    .keyStatus_20_valid       (debounce_1_keyStatus_20_valid     ), //o
    .keyStatus_20_payload     (debounce_1_keyStatus_20_payload   ), //o
    .keyStatus_21_valid       (debounce_1_keyStatus_21_valid     ), //o
    .keyStatus_21_payload     (debounce_1_keyStatus_21_payload   ), //o
    .keyStatus_22_valid       (debounce_1_keyStatus_22_valid     ), //o
    .keyStatus_22_payload     (debounce_1_keyStatus_22_payload   ), //o
    .keyStatus_23_valid       (debounce_1_keyStatus_23_valid     ), //o
    .keyStatus_23_payload     (debounce_1_keyStatus_23_payload   ), //o
    .keyStatus_24_valid       (debounce_1_keyStatus_24_valid     ), //o
    .keyStatus_24_payload     (debounce_1_keyStatus_24_payload   ), //o
    .keyStatus_25_valid       (debounce_1_keyStatus_25_valid     ), //o
    .keyStatus_25_payload     (debounce_1_keyStatus_25_payload   ), //o
    .keyStatus_26_valid       (debounce_1_keyStatus_26_valid     ), //o
    .keyStatus_26_payload     (debounce_1_keyStatus_26_payload   ), //o
    .keyStatus_27_valid       (debounce_1_keyStatus_27_valid     ), //o
    .keyStatus_27_payload     (debounce_1_keyStatus_27_payload   ), //o
    .keyStatus_28_valid       (debounce_1_keyStatus_28_valid     ), //o
    .keyStatus_28_payload     (debounce_1_keyStatus_28_payload   ), //o
    .keyStatus_29_valid       (debounce_1_keyStatus_29_valid     ), //o
    .keyStatus_29_payload     (debounce_1_keyStatus_29_payload   ), //o
    .keyStatus_30_valid       (debounce_1_keyStatus_30_valid     ), //o
    .keyStatus_30_payload     (debounce_1_keyStatus_30_payload   ), //o
    .keyStatus_31_valid       (debounce_1_keyStatus_31_valid     ), //o
    .keyStatus_31_payload     (debounce_1_keyStatus_31_payload   ), //o
    .keyStatus_32_valid       (debounce_1_keyStatus_32_valid     ), //o
    .keyStatus_32_payload     (debounce_1_keyStatus_32_payload   ), //o
    .keyStatus_33_valid       (debounce_1_keyStatus_33_valid     ), //o
    .keyStatus_33_payload     (debounce_1_keyStatus_33_payload   ), //o
    .keyStatus_34_valid       (debounce_1_keyStatus_34_valid     ), //o
    .keyStatus_34_payload     (debounce_1_keyStatus_34_payload   ), //o
    .keyStatus_35_valid       (debounce_1_keyStatus_35_valid     ), //o
    .keyStatus_35_payload     (debounce_1_keyStatus_35_payload   ), //o
    .keyStatus_36_valid       (debounce_1_keyStatus_36_valid     ), //o
    .keyStatus_36_payload     (debounce_1_keyStatus_36_payload   ), //o
    .keyStatus_37_valid       (debounce_1_keyStatus_37_valid     ), //o
    .keyStatus_37_payload     (debounce_1_keyStatus_37_payload   ), //o
    .keyStatus_38_valid       (debounce_1_keyStatus_38_valid     ), //o
    .keyStatus_38_payload     (debounce_1_keyStatus_38_payload   ), //o
    .keyStatus_39_valid       (debounce_1_keyStatus_39_valid     ), //o
    .keyStatus_39_payload     (debounce_1_keyStatus_39_payload   ), //o
    .keyStatus_40_valid       (debounce_1_keyStatus_40_valid     ), //o
    .keyStatus_40_payload     (debounce_1_keyStatus_40_payload   ), //o
    .keyStatus_41_valid       (debounce_1_keyStatus_41_valid     ), //o
    .keyStatus_41_payload     (debounce_1_keyStatus_41_payload   ), //o
    .keyStatus_42_valid       (debounce_1_keyStatus_42_valid     ), //o
    .keyStatus_42_payload     (debounce_1_keyStatus_42_payload   ), //o
    .keyStatus_43_valid       (debounce_1_keyStatus_43_valid     ), //o
    .keyStatus_43_payload     (debounce_1_keyStatus_43_payload   ), //o
    .keyStatus_44_valid       (debounce_1_keyStatus_44_valid     ), //o
    .keyStatus_44_payload     (debounce_1_keyStatus_44_payload   ), //o
    .keyStatus_45_valid       (debounce_1_keyStatus_45_valid     ), //o
    .keyStatus_45_payload     (debounce_1_keyStatus_45_payload   ), //o
    .keyStatus_46_valid       (debounce_1_keyStatus_46_valid     ), //o
    .keyStatus_46_payload     (debounce_1_keyStatus_46_payload   ), //o
    .keyStatus_47_valid       (debounce_1_keyStatus_47_valid     ), //o
    .keyStatus_47_payload     (debounce_1_keyStatus_47_payload   ), //o
    .keyStatus_48_valid       (debounce_1_keyStatus_48_valid     ), //o
    .keyStatus_48_payload     (debounce_1_keyStatus_48_payload   ), //o
    .keyStatus_49_valid       (debounce_1_keyStatus_49_valid     ), //o
    .keyStatus_49_payload     (debounce_1_keyStatus_49_payload   ), //o
    .keyStatus_50_valid       (debounce_1_keyStatus_50_valid     ), //o
    .keyStatus_50_payload     (debounce_1_keyStatus_50_payload   ), //o
    .keyStatus_51_valid       (debounce_1_keyStatus_51_valid     ), //o
    .keyStatus_51_payload     (debounce_1_keyStatus_51_payload   ), //o
    .keyStatus_52_valid       (debounce_1_keyStatus_52_valid     ), //o
    .keyStatus_52_payload     (debounce_1_keyStatus_52_payload   ), //o
    .keyStatus_53_valid       (debounce_1_keyStatus_53_valid     ), //o
    .keyStatus_53_payload     (debounce_1_keyStatus_53_payload   ), //o
    .keyStatus_54_valid       (debounce_1_keyStatus_54_valid     ), //o
    .keyStatus_54_payload     (debounce_1_keyStatus_54_payload   ), //o
    .keyStatus_55_valid       (debounce_1_keyStatus_55_valid     ), //o
    .keyStatus_55_payload     (debounce_1_keyStatus_55_payload   ), //o
    .keyStatus_56_valid       (debounce_1_keyStatus_56_valid     ), //o
    .keyStatus_56_payload     (debounce_1_keyStatus_56_payload   ), //o
    .keyStatus_57_valid       (debounce_1_keyStatus_57_valid     ), //o
    .keyStatus_57_payload     (debounce_1_keyStatus_57_payload   ), //o
    .keyStatus_58_valid       (debounce_1_keyStatus_58_valid     ), //o
    .keyStatus_58_payload     (debounce_1_keyStatus_58_payload   ), //o
    .keyStatus_59_valid       (debounce_1_keyStatus_59_valid     ), //o
    .keyStatus_59_payload     (debounce_1_keyStatus_59_payload   ), //o
    .keyStatus_60_valid       (debounce_1_keyStatus_60_valid     ), //o
    .keyStatus_60_payload     (debounce_1_keyStatus_60_payload   ), //o
    .keyStatus_61_valid       (debounce_1_keyStatus_61_valid     ), //o
    .keyStatus_61_payload     (debounce_1_keyStatus_61_payload   ), //o
    .keyStatus_62_valid       (debounce_1_keyStatus_62_valid     ), //o
    .keyStatus_62_payload     (debounce_1_keyStatus_62_payload   ), //o
    .keyStatus_63_valid       (debounce_1_keyStatus_63_valid     ), //o
    .keyStatus_63_payload     (debounce_1_keyStatus_63_payload   ), //o
    .keyStatus_64_valid       (debounce_1_keyStatus_64_valid     ), //o
    .keyStatus_64_payload     (debounce_1_keyStatus_64_payload   ), //o
    .keyStatus_65_valid       (debounce_1_keyStatus_65_valid     ), //o
    .keyStatus_65_payload     (debounce_1_keyStatus_65_payload   ), //o
    .keyStatus_66_valid       (debounce_1_keyStatus_66_valid     ), //o
    .keyStatus_66_payload     (debounce_1_keyStatus_66_payload   ), //o
    .keyStatus_67_valid       (debounce_1_keyStatus_67_valid     ), //o
    .keyStatus_67_payload     (debounce_1_keyStatus_67_payload   ), //o
    .keyStatus_68_valid       (debounce_1_keyStatus_68_valid     ), //o
    .keyStatus_68_payload     (debounce_1_keyStatus_68_payload   ), //o
    .keyStatus_69_valid       (debounce_1_keyStatus_69_valid     ), //o
    .keyStatus_69_payload     (debounce_1_keyStatus_69_payload   ), //o
    .keyStatus_70_valid       (debounce_1_keyStatus_70_valid     ), //o
    .keyStatus_70_payload     (debounce_1_keyStatus_70_payload   ), //o
    .keyStatus_71_valid       (debounce_1_keyStatus_71_valid     ), //o
    .keyStatus_71_payload     (debounce_1_keyStatus_71_payload   ), //o
    .keyStatus_72_valid       (debounce_1_keyStatus_72_valid     ), //o
    .keyStatus_72_payload     (debounce_1_keyStatus_72_payload   ), //o
    .keyStatus_73_valid       (debounce_1_keyStatus_73_valid     ), //o
    .keyStatus_73_payload     (debounce_1_keyStatus_73_payload   ), //o
    .keyStatus_74_valid       (debounce_1_keyStatus_74_valid     ), //o
    .keyStatus_74_payload     (debounce_1_keyStatus_74_payload   ), //o
    .keyStatus_75_valid       (debounce_1_keyStatus_75_valid     ), //o
    .keyStatus_75_payload     (debounce_1_keyStatus_75_payload   ), //o
    .keyStatus_76_valid       (debounce_1_keyStatus_76_valid     ), //o
    .keyStatus_76_payload     (debounce_1_keyStatus_76_payload   ), //o
    .keyStatus_77_valid       (debounce_1_keyStatus_77_valid     ), //o
    .keyStatus_77_payload     (debounce_1_keyStatus_77_payload   ), //o
    .keyStatus_78_valid       (debounce_1_keyStatus_78_valid     ), //o
    .keyStatus_78_payload     (debounce_1_keyStatus_78_payload   ), //o
    .keyStatus_79_valid       (debounce_1_keyStatus_79_valid     ), //o
    .keyStatus_79_payload     (debounce_1_keyStatus_79_payload   ), //o
    .keyStatus_80_valid       (debounce_1_keyStatus_80_valid     ), //o
    .keyStatus_80_payload     (debounce_1_keyStatus_80_payload   ), //o
    .keyStatus_81_valid       (debounce_1_keyStatus_81_valid     ), //o
    .keyStatus_81_payload     (debounce_1_keyStatus_81_payload   ), //o
    .keyStatus_82_valid       (debounce_1_keyStatus_82_valid     ), //o
    .keyStatus_82_payload     (debounce_1_keyStatus_82_payload   ), //o
    .keyStatus_83_valid       (debounce_1_keyStatus_83_valid     ), //o
    .keyStatus_83_payload     (debounce_1_keyStatus_83_payload   ), //o
    .keyStatus_84_valid       (debounce_1_keyStatus_84_valid     ), //o
    .keyStatus_84_payload     (debounce_1_keyStatus_84_payload   ), //o
    .keyStatus_85_valid       (debounce_1_keyStatus_85_valid     ), //o
    .keyStatus_85_payload     (debounce_1_keyStatus_85_payload   ), //o
    .keyStatus_86_valid       (debounce_1_keyStatus_86_valid     ), //o
    .keyStatus_86_payload     (debounce_1_keyStatus_86_payload   ), //o
    .keyStatus_87_valid       (debounce_1_keyStatus_87_valid     ), //o
    .keyStatus_87_payload     (debounce_1_keyStatus_87_payload   ), //o
    .keyStatus_88_valid       (debounce_1_keyStatus_88_valid     ), //o
    .keyStatus_88_payload     (debounce_1_keyStatus_88_payload   ), //o
    .keyStatus_89_valid       (debounce_1_keyStatus_89_valid     ), //o
    .keyStatus_89_payload     (debounce_1_keyStatus_89_payload   ), //o
    .keyStatus_90_valid       (debounce_1_keyStatus_90_valid     ), //o
    .keyStatus_90_payload     (debounce_1_keyStatus_90_payload   ), //o
    .keyStatus_91_valid       (debounce_1_keyStatus_91_valid     ), //o
    .keyStatus_91_payload     (debounce_1_keyStatus_91_payload   ), //o
    .keyStatus_92_valid       (debounce_1_keyStatus_92_valid     ), //o
    .keyStatus_92_payload     (debounce_1_keyStatus_92_payload   ), //o
    .keyStatus_93_valid       (debounce_1_keyStatus_93_valid     ), //o
    .keyStatus_93_payload     (debounce_1_keyStatus_93_payload   ), //o
    .keyStatus_94_valid       (debounce_1_keyStatus_94_valid     ), //o
    .keyStatus_94_payload     (debounce_1_keyStatus_94_payload   ), //o
    .keyStatus_95_valid       (debounce_1_keyStatus_95_valid     ), //o
    .keyStatus_95_payload     (debounce_1_keyStatus_95_payload   ), //o
    .keyStatus_96_valid       (debounce_1_keyStatus_96_valid     ), //o
    .keyStatus_96_payload     (debounce_1_keyStatus_96_payload   ), //o
    .keyStatus_97_valid       (debounce_1_keyStatus_97_valid     ), //o
    .keyStatus_97_payload     (debounce_1_keyStatus_97_payload   ), //o
    .keyStatus_98_valid       (debounce_1_keyStatus_98_valid     ), //o
    .keyStatus_98_payload     (debounce_1_keyStatus_98_payload   ), //o
    .keyStatus_99_valid       (debounce_1_keyStatus_99_valid     ), //o
    .keyStatus_99_payload     (debounce_1_keyStatus_99_payload   ), //o
    .keyStatus_100_valid      (debounce_1_keyStatus_100_valid    ), //o
    .keyStatus_100_payload    (debounce_1_keyStatus_100_payload  ), //o
    .keyStatus_101_valid      (debounce_1_keyStatus_101_valid    ), //o
    .keyStatus_101_payload    (debounce_1_keyStatus_101_payload  ), //o
    .keyStatus_102_valid      (debounce_1_keyStatus_102_valid    ), //o
    .keyStatus_102_payload    (debounce_1_keyStatus_102_payload  ), //o
    .CLK_50                   (CLK_50                            ), //i
    ._zz_3                    (_zz_1                             )  //i
  );
  always @(*) begin
    case(_zz_6)
      7'b0000000 : begin
        _zz_9 = keyStatus_0_valid;
        _zz_10 = keyStatus_0_payload;
      end
      7'b0000001 : begin
        _zz_9 = keyStatus_1_valid;
        _zz_10 = keyStatus_1_payload;
      end
      7'b0000010 : begin
        _zz_9 = keyStatus_2_valid;
        _zz_10 = keyStatus_2_payload;
      end
      7'b0000011 : begin
        _zz_9 = keyStatus_3_valid;
        _zz_10 = keyStatus_3_payload;
      end
      7'b0000100 : begin
        _zz_9 = keyStatus_4_valid;
        _zz_10 = keyStatus_4_payload;
      end
      7'b0000101 : begin
        _zz_9 = keyStatus_5_valid;
        _zz_10 = keyStatus_5_payload;
      end
      7'b0000110 : begin
        _zz_9 = keyStatus_6_valid;
        _zz_10 = keyStatus_6_payload;
      end
      7'b0000111 : begin
        _zz_9 = keyStatus_7_valid;
        _zz_10 = keyStatus_7_payload;
      end
      7'b0001000 : begin
        _zz_9 = keyStatus_8_valid;
        _zz_10 = keyStatus_8_payload;
      end
      7'b0001001 : begin
        _zz_9 = keyStatus_9_valid;
        _zz_10 = keyStatus_9_payload;
      end
      7'b0001010 : begin
        _zz_9 = keyStatus_10_valid;
        _zz_10 = keyStatus_10_payload;
      end
      7'b0001011 : begin
        _zz_9 = keyStatus_11_valid;
        _zz_10 = keyStatus_11_payload;
      end
      7'b0001100 : begin
        _zz_9 = keyStatus_12_valid;
        _zz_10 = keyStatus_12_payload;
      end
      7'b0001101 : begin
        _zz_9 = keyStatus_13_valid;
        _zz_10 = keyStatus_13_payload;
      end
      7'b0001110 : begin
        _zz_9 = keyStatus_14_valid;
        _zz_10 = keyStatus_14_payload;
      end
      7'b0001111 : begin
        _zz_9 = keyStatus_15_valid;
        _zz_10 = keyStatus_15_payload;
      end
      7'b0010000 : begin
        _zz_9 = keyStatus_16_valid;
        _zz_10 = keyStatus_16_payload;
      end
      7'b0010001 : begin
        _zz_9 = keyStatus_17_valid;
        _zz_10 = keyStatus_17_payload;
      end
      7'b0010010 : begin
        _zz_9 = keyStatus_18_valid;
        _zz_10 = keyStatus_18_payload;
      end
      7'b0010011 : begin
        _zz_9 = keyStatus_19_valid;
        _zz_10 = keyStatus_19_payload;
      end
      7'b0010100 : begin
        _zz_9 = keyStatus_20_valid;
        _zz_10 = keyStatus_20_payload;
      end
      7'b0010101 : begin
        _zz_9 = keyStatus_21_valid;
        _zz_10 = keyStatus_21_payload;
      end
      7'b0010110 : begin
        _zz_9 = keyStatus_22_valid;
        _zz_10 = keyStatus_22_payload;
      end
      7'b0010111 : begin
        _zz_9 = keyStatus_23_valid;
        _zz_10 = keyStatus_23_payload;
      end
      7'b0011000 : begin
        _zz_9 = keyStatus_24_valid;
        _zz_10 = keyStatus_24_payload;
      end
      7'b0011001 : begin
        _zz_9 = keyStatus_25_valid;
        _zz_10 = keyStatus_25_payload;
      end
      7'b0011010 : begin
        _zz_9 = keyStatus_26_valid;
        _zz_10 = keyStatus_26_payload;
      end
      7'b0011011 : begin
        _zz_9 = keyStatus_27_valid;
        _zz_10 = keyStatus_27_payload;
      end
      7'b0011100 : begin
        _zz_9 = keyStatus_28_valid;
        _zz_10 = keyStatus_28_payload;
      end
      7'b0011101 : begin
        _zz_9 = keyStatus_29_valid;
        _zz_10 = keyStatus_29_payload;
      end
      7'b0011110 : begin
        _zz_9 = keyStatus_30_valid;
        _zz_10 = keyStatus_30_payload;
      end
      7'b0011111 : begin
        _zz_9 = keyStatus_31_valid;
        _zz_10 = keyStatus_31_payload;
      end
      7'b0100000 : begin
        _zz_9 = keyStatus_32_valid;
        _zz_10 = keyStatus_32_payload;
      end
      7'b0100001 : begin
        _zz_9 = keyStatus_33_valid;
        _zz_10 = keyStatus_33_payload;
      end
      7'b0100010 : begin
        _zz_9 = keyStatus_34_valid;
        _zz_10 = keyStatus_34_payload;
      end
      7'b0100011 : begin
        _zz_9 = keyStatus_35_valid;
        _zz_10 = keyStatus_35_payload;
      end
      7'b0100100 : begin
        _zz_9 = keyStatus_36_valid;
        _zz_10 = keyStatus_36_payload;
      end
      7'b0100101 : begin
        _zz_9 = keyStatus_37_valid;
        _zz_10 = keyStatus_37_payload;
      end
      7'b0100110 : begin
        _zz_9 = keyStatus_38_valid;
        _zz_10 = keyStatus_38_payload;
      end
      7'b0100111 : begin
        _zz_9 = keyStatus_39_valid;
        _zz_10 = keyStatus_39_payload;
      end
      7'b0101000 : begin
        _zz_9 = keyStatus_40_valid;
        _zz_10 = keyStatus_40_payload;
      end
      7'b0101001 : begin
        _zz_9 = keyStatus_41_valid;
        _zz_10 = keyStatus_41_payload;
      end
      7'b0101010 : begin
        _zz_9 = keyStatus_42_valid;
        _zz_10 = keyStatus_42_payload;
      end
      7'b0101011 : begin
        _zz_9 = keyStatus_43_valid;
        _zz_10 = keyStatus_43_payload;
      end
      7'b0101100 : begin
        _zz_9 = keyStatus_44_valid;
        _zz_10 = keyStatus_44_payload;
      end
      7'b0101101 : begin
        _zz_9 = keyStatus_45_valid;
        _zz_10 = keyStatus_45_payload;
      end
      7'b0101110 : begin
        _zz_9 = keyStatus_46_valid;
        _zz_10 = keyStatus_46_payload;
      end
      7'b0101111 : begin
        _zz_9 = keyStatus_47_valid;
        _zz_10 = keyStatus_47_payload;
      end
      7'b0110000 : begin
        _zz_9 = keyStatus_48_valid;
        _zz_10 = keyStatus_48_payload;
      end
      7'b0110001 : begin
        _zz_9 = keyStatus_49_valid;
        _zz_10 = keyStatus_49_payload;
      end
      7'b0110010 : begin
        _zz_9 = keyStatus_50_valid;
        _zz_10 = keyStatus_50_payload;
      end
      7'b0110011 : begin
        _zz_9 = keyStatus_51_valid;
        _zz_10 = keyStatus_51_payload;
      end
      7'b0110100 : begin
        _zz_9 = keyStatus_52_valid;
        _zz_10 = keyStatus_52_payload;
      end
      7'b0110101 : begin
        _zz_9 = keyStatus_53_valid;
        _zz_10 = keyStatus_53_payload;
      end
      7'b0110110 : begin
        _zz_9 = keyStatus_54_valid;
        _zz_10 = keyStatus_54_payload;
      end
      7'b0110111 : begin
        _zz_9 = keyStatus_55_valid;
        _zz_10 = keyStatus_55_payload;
      end
      7'b0111000 : begin
        _zz_9 = keyStatus_56_valid;
        _zz_10 = keyStatus_56_payload;
      end
      7'b0111001 : begin
        _zz_9 = keyStatus_57_valid;
        _zz_10 = keyStatus_57_payload;
      end
      7'b0111010 : begin
        _zz_9 = keyStatus_58_valid;
        _zz_10 = keyStatus_58_payload;
      end
      7'b0111011 : begin
        _zz_9 = keyStatus_59_valid;
        _zz_10 = keyStatus_59_payload;
      end
      7'b0111100 : begin
        _zz_9 = keyStatus_60_valid;
        _zz_10 = keyStatus_60_payload;
      end
      7'b0111101 : begin
        _zz_9 = keyStatus_61_valid;
        _zz_10 = keyStatus_61_payload;
      end
      7'b0111110 : begin
        _zz_9 = keyStatus_62_valid;
        _zz_10 = keyStatus_62_payload;
      end
      7'b0111111 : begin
        _zz_9 = keyStatus_63_valid;
        _zz_10 = keyStatus_63_payload;
      end
      7'b1000000 : begin
        _zz_9 = keyStatus_64_valid;
        _zz_10 = keyStatus_64_payload;
      end
      7'b1000001 : begin
        _zz_9 = keyStatus_65_valid;
        _zz_10 = keyStatus_65_payload;
      end
      7'b1000010 : begin
        _zz_9 = keyStatus_66_valid;
        _zz_10 = keyStatus_66_payload;
      end
      7'b1000011 : begin
        _zz_9 = keyStatus_67_valid;
        _zz_10 = keyStatus_67_payload;
      end
      7'b1000100 : begin
        _zz_9 = keyStatus_68_valid;
        _zz_10 = keyStatus_68_payload;
      end
      7'b1000101 : begin
        _zz_9 = keyStatus_69_valid;
        _zz_10 = keyStatus_69_payload;
      end
      7'b1000110 : begin
        _zz_9 = keyStatus_70_valid;
        _zz_10 = keyStatus_70_payload;
      end
      7'b1000111 : begin
        _zz_9 = keyStatus_71_valid;
        _zz_10 = keyStatus_71_payload;
      end
      7'b1001000 : begin
        _zz_9 = keyStatus_72_valid;
        _zz_10 = keyStatus_72_payload;
      end
      7'b1001001 : begin
        _zz_9 = keyStatus_73_valid;
        _zz_10 = keyStatus_73_payload;
      end
      7'b1001010 : begin
        _zz_9 = keyStatus_74_valid;
        _zz_10 = keyStatus_74_payload;
      end
      7'b1001011 : begin
        _zz_9 = keyStatus_75_valid;
        _zz_10 = keyStatus_75_payload;
      end
      7'b1001100 : begin
        _zz_9 = keyStatus_76_valid;
        _zz_10 = keyStatus_76_payload;
      end
      7'b1001101 : begin
        _zz_9 = keyStatus_77_valid;
        _zz_10 = keyStatus_77_payload;
      end
      7'b1001110 : begin
        _zz_9 = keyStatus_78_valid;
        _zz_10 = keyStatus_78_payload;
      end
      7'b1001111 : begin
        _zz_9 = keyStatus_79_valid;
        _zz_10 = keyStatus_79_payload;
      end
      7'b1010000 : begin
        _zz_9 = keyStatus_80_valid;
        _zz_10 = keyStatus_80_payload;
      end
      7'b1010001 : begin
        _zz_9 = keyStatus_81_valid;
        _zz_10 = keyStatus_81_payload;
      end
      7'b1010010 : begin
        _zz_9 = keyStatus_82_valid;
        _zz_10 = keyStatus_82_payload;
      end
      7'b1010011 : begin
        _zz_9 = keyStatus_83_valid;
        _zz_10 = keyStatus_83_payload;
      end
      7'b1010100 : begin
        _zz_9 = keyStatus_84_valid;
        _zz_10 = keyStatus_84_payload;
      end
      7'b1010101 : begin
        _zz_9 = keyStatus_85_valid;
        _zz_10 = keyStatus_85_payload;
      end
      7'b1010110 : begin
        _zz_9 = keyStatus_86_valid;
        _zz_10 = keyStatus_86_payload;
      end
      7'b1010111 : begin
        _zz_9 = keyStatus_87_valid;
        _zz_10 = keyStatus_87_payload;
      end
      7'b1011000 : begin
        _zz_9 = keyStatus_88_valid;
        _zz_10 = keyStatus_88_payload;
      end
      7'b1011001 : begin
        _zz_9 = keyStatus_89_valid;
        _zz_10 = keyStatus_89_payload;
      end
      7'b1011010 : begin
        _zz_9 = keyStatus_90_valid;
        _zz_10 = keyStatus_90_payload;
      end
      7'b1011011 : begin
        _zz_9 = keyStatus_91_valid;
        _zz_10 = keyStatus_91_payload;
      end
      7'b1011100 : begin
        _zz_9 = keyStatus_92_valid;
        _zz_10 = keyStatus_92_payload;
      end
      7'b1011101 : begin
        _zz_9 = keyStatus_93_valid;
        _zz_10 = keyStatus_93_payload;
      end
      7'b1011110 : begin
        _zz_9 = keyStatus_94_valid;
        _zz_10 = keyStatus_94_payload;
      end
      7'b1011111 : begin
        _zz_9 = keyStatus_95_valid;
        _zz_10 = keyStatus_95_payload;
      end
      7'b1100000 : begin
        _zz_9 = keyStatus_96_valid;
        _zz_10 = keyStatus_96_payload;
      end
      7'b1100001 : begin
        _zz_9 = keyStatus_97_valid;
        _zz_10 = keyStatus_97_payload;
      end
      7'b1100010 : begin
        _zz_9 = keyStatus_98_valid;
        _zz_10 = keyStatus_98_payload;
      end
      7'b1100011 : begin
        _zz_9 = keyStatus_99_valid;
        _zz_10 = keyStatus_99_payload;
      end
      7'b1100100 : begin
        _zz_9 = keyStatus_100_valid;
        _zz_10 = keyStatus_100_payload;
      end
      7'b1100101 : begin
        _zz_9 = keyStatus_101_valid;
        _zz_10 = keyStatus_101_payload;
      end
      default : begin
        _zz_9 = keyStatus_102_valid;
        _zz_10 = keyStatus_102_payload;
      end
    endcase
  end

  assign keyBits = {{keyStatus_102_payload,keyStatus_102_valid},{{keyStatus_101_payload,keyStatus_101_valid},{{keyStatus_100_payload,keyStatus_100_valid},{{keyStatus_99_payload,keyStatus_99_valid},{{keyStatus_98_payload,keyStatus_98_valid},{{_zz_15,_zz_16},{_zz_17,_zz_18}}}}}}};
  always @ (*) begin
    clkScan_stateRise = 1'b0;
    if(clkScan_counter_willOverflow)begin
      clkScan_stateRise = (! clkScan_state);
    end
    if(clkScan_state)begin
      clkScan_stateRise = 1'b0;
    end
  end

  always @ (*) begin
    clkScan_counter_willClear = 1'b0;
    if(clkScan_state)begin
      clkScan_counter_willClear = 1'b1;
    end
  end

  assign clkScan_counter_willOverflowIfInc = (clkScan_counter_value == 11'h681);
  assign clkScan_counter_willOverflow = (clkScan_counter_willOverflowIfInc && clkScan_counter_willIncrement);
  always @ (*) begin
    if(clkScan_counter_willOverflow)begin
      clkScan_counter_valueNext = 11'h0;
    end else begin
      clkScan_counter_valueNext = (clkScan_counter_value + _zz_12);
    end
    if(clkScan_counter_willClear)begin
      clkScan_counter_valueNext = 11'h0;
    end
  end

  assign clkScan_counter_willIncrement = 1'b1;
  assign ROW = scanK_ROW;
  assign keyStatus_0_valid = debounce_1_keyStatus_0_valid;
  assign keyStatus_0_payload = debounce_1_keyStatus_0_payload;
  assign keyStatus_1_valid = debounce_1_keyStatus_1_valid;
  assign keyStatus_1_payload = debounce_1_keyStatus_1_payload;
  assign keyStatus_2_valid = debounce_1_keyStatus_2_valid;
  assign keyStatus_2_payload = debounce_1_keyStatus_2_payload;
  assign keyStatus_3_valid = debounce_1_keyStatus_3_valid;
  assign keyStatus_3_payload = debounce_1_keyStatus_3_payload;
  assign keyStatus_4_valid = debounce_1_keyStatus_4_valid;
  assign keyStatus_4_payload = debounce_1_keyStatus_4_payload;
  assign keyStatus_5_valid = debounce_1_keyStatus_5_valid;
  assign keyStatus_5_payload = debounce_1_keyStatus_5_payload;
  assign keyStatus_6_valid = debounce_1_keyStatus_6_valid;
  assign keyStatus_6_payload = debounce_1_keyStatus_6_payload;
  assign keyStatus_7_valid = debounce_1_keyStatus_7_valid;
  assign keyStatus_7_payload = debounce_1_keyStatus_7_payload;
  assign keyStatus_8_valid = debounce_1_keyStatus_8_valid;
  assign keyStatus_8_payload = debounce_1_keyStatus_8_payload;
  assign keyStatus_9_valid = debounce_1_keyStatus_9_valid;
  assign keyStatus_9_payload = debounce_1_keyStatus_9_payload;
  assign keyStatus_10_valid = debounce_1_keyStatus_10_valid;
  assign keyStatus_10_payload = debounce_1_keyStatus_10_payload;
  assign keyStatus_11_valid = debounce_1_keyStatus_11_valid;
  assign keyStatus_11_payload = debounce_1_keyStatus_11_payload;
  assign keyStatus_12_valid = debounce_1_keyStatus_12_valid;
  assign keyStatus_12_payload = debounce_1_keyStatus_12_payload;
  assign keyStatus_13_valid = debounce_1_keyStatus_13_valid;
  assign keyStatus_13_payload = debounce_1_keyStatus_13_payload;
  assign keyStatus_14_valid = debounce_1_keyStatus_14_valid;
  assign keyStatus_14_payload = debounce_1_keyStatus_14_payload;
  assign keyStatus_15_valid = debounce_1_keyStatus_15_valid;
  assign keyStatus_15_payload = debounce_1_keyStatus_15_payload;
  assign keyStatus_16_valid = debounce_1_keyStatus_16_valid;
  assign keyStatus_16_payload = debounce_1_keyStatus_16_payload;
  assign keyStatus_17_valid = debounce_1_keyStatus_17_valid;
  assign keyStatus_17_payload = debounce_1_keyStatus_17_payload;
  assign keyStatus_18_valid = debounce_1_keyStatus_18_valid;
  assign keyStatus_18_payload = debounce_1_keyStatus_18_payload;
  assign keyStatus_19_valid = debounce_1_keyStatus_19_valid;
  assign keyStatus_19_payload = debounce_1_keyStatus_19_payload;
  assign keyStatus_20_valid = debounce_1_keyStatus_20_valid;
  assign keyStatus_20_payload = debounce_1_keyStatus_20_payload;
  assign keyStatus_21_valid = debounce_1_keyStatus_21_valid;
  assign keyStatus_21_payload = debounce_1_keyStatus_21_payload;
  assign keyStatus_22_valid = debounce_1_keyStatus_22_valid;
  assign keyStatus_22_payload = debounce_1_keyStatus_22_payload;
  assign keyStatus_23_valid = debounce_1_keyStatus_23_valid;
  assign keyStatus_23_payload = debounce_1_keyStatus_23_payload;
  assign keyStatus_24_valid = debounce_1_keyStatus_24_valid;
  assign keyStatus_24_payload = debounce_1_keyStatus_24_payload;
  assign keyStatus_25_valid = debounce_1_keyStatus_25_valid;
  assign keyStatus_25_payload = debounce_1_keyStatus_25_payload;
  assign keyStatus_26_valid = debounce_1_keyStatus_26_valid;
  assign keyStatus_26_payload = debounce_1_keyStatus_26_payload;
  assign keyStatus_27_valid = debounce_1_keyStatus_27_valid;
  assign keyStatus_27_payload = debounce_1_keyStatus_27_payload;
  assign keyStatus_28_valid = debounce_1_keyStatus_28_valid;
  assign keyStatus_28_payload = debounce_1_keyStatus_28_payload;
  assign keyStatus_29_valid = debounce_1_keyStatus_29_valid;
  assign keyStatus_29_payload = debounce_1_keyStatus_29_payload;
  assign keyStatus_30_valid = debounce_1_keyStatus_30_valid;
  assign keyStatus_30_payload = debounce_1_keyStatus_30_payload;
  assign keyStatus_31_valid = debounce_1_keyStatus_31_valid;
  assign keyStatus_31_payload = debounce_1_keyStatus_31_payload;
  assign keyStatus_32_valid = debounce_1_keyStatus_32_valid;
  assign keyStatus_32_payload = debounce_1_keyStatus_32_payload;
  assign keyStatus_33_valid = debounce_1_keyStatus_33_valid;
  assign keyStatus_33_payload = debounce_1_keyStatus_33_payload;
  assign keyStatus_34_valid = debounce_1_keyStatus_34_valid;
  assign keyStatus_34_payload = debounce_1_keyStatus_34_payload;
  assign keyStatus_35_valid = debounce_1_keyStatus_35_valid;
  assign keyStatus_35_payload = debounce_1_keyStatus_35_payload;
  assign keyStatus_36_valid = debounce_1_keyStatus_36_valid;
  assign keyStatus_36_payload = debounce_1_keyStatus_36_payload;
  assign keyStatus_37_valid = debounce_1_keyStatus_37_valid;
  assign keyStatus_37_payload = debounce_1_keyStatus_37_payload;
  assign keyStatus_38_valid = debounce_1_keyStatus_38_valid;
  assign keyStatus_38_payload = debounce_1_keyStatus_38_payload;
  assign keyStatus_39_valid = debounce_1_keyStatus_39_valid;
  assign keyStatus_39_payload = debounce_1_keyStatus_39_payload;
  assign keyStatus_40_valid = debounce_1_keyStatus_40_valid;
  assign keyStatus_40_payload = debounce_1_keyStatus_40_payload;
  assign keyStatus_41_valid = debounce_1_keyStatus_41_valid;
  assign keyStatus_41_payload = debounce_1_keyStatus_41_payload;
  assign keyStatus_42_valid = debounce_1_keyStatus_42_valid;
  assign keyStatus_42_payload = debounce_1_keyStatus_42_payload;
  assign keyStatus_43_valid = debounce_1_keyStatus_43_valid;
  assign keyStatus_43_payload = debounce_1_keyStatus_43_payload;
  assign keyStatus_44_valid = debounce_1_keyStatus_44_valid;
  assign keyStatus_44_payload = debounce_1_keyStatus_44_payload;
  assign keyStatus_45_valid = debounce_1_keyStatus_45_valid;
  assign keyStatus_45_payload = debounce_1_keyStatus_45_payload;
  assign keyStatus_46_valid = debounce_1_keyStatus_46_valid;
  assign keyStatus_46_payload = debounce_1_keyStatus_46_payload;
  assign keyStatus_47_valid = debounce_1_keyStatus_47_valid;
  assign keyStatus_47_payload = debounce_1_keyStatus_47_payload;
  assign keyStatus_48_valid = debounce_1_keyStatus_48_valid;
  assign keyStatus_48_payload = debounce_1_keyStatus_48_payload;
  assign keyStatus_49_valid = debounce_1_keyStatus_49_valid;
  assign keyStatus_49_payload = debounce_1_keyStatus_49_payload;
  assign keyStatus_50_valid = debounce_1_keyStatus_50_valid;
  assign keyStatus_50_payload = debounce_1_keyStatus_50_payload;
  assign keyStatus_51_valid = debounce_1_keyStatus_51_valid;
  assign keyStatus_51_payload = debounce_1_keyStatus_51_payload;
  assign keyStatus_52_valid = debounce_1_keyStatus_52_valid;
  assign keyStatus_52_payload = debounce_1_keyStatus_52_payload;
  assign keyStatus_53_valid = debounce_1_keyStatus_53_valid;
  assign keyStatus_53_payload = debounce_1_keyStatus_53_payload;
  assign keyStatus_54_valid = debounce_1_keyStatus_54_valid;
  assign keyStatus_54_payload = debounce_1_keyStatus_54_payload;
  assign keyStatus_55_valid = debounce_1_keyStatus_55_valid;
  assign keyStatus_55_payload = debounce_1_keyStatus_55_payload;
  assign keyStatus_56_valid = debounce_1_keyStatus_56_valid;
  assign keyStatus_56_payload = debounce_1_keyStatus_56_payload;
  assign keyStatus_57_valid = debounce_1_keyStatus_57_valid;
  assign keyStatus_57_payload = debounce_1_keyStatus_57_payload;
  assign keyStatus_58_valid = debounce_1_keyStatus_58_valid;
  assign keyStatus_58_payload = debounce_1_keyStatus_58_payload;
  assign keyStatus_59_valid = debounce_1_keyStatus_59_valid;
  assign keyStatus_59_payload = debounce_1_keyStatus_59_payload;
  assign keyStatus_60_valid = debounce_1_keyStatus_60_valid;
  assign keyStatus_60_payload = debounce_1_keyStatus_60_payload;
  assign keyStatus_61_valid = debounce_1_keyStatus_61_valid;
  assign keyStatus_61_payload = debounce_1_keyStatus_61_payload;
  assign keyStatus_62_valid = debounce_1_keyStatus_62_valid;
  assign keyStatus_62_payload = debounce_1_keyStatus_62_payload;
  assign keyStatus_63_valid = debounce_1_keyStatus_63_valid;
  assign keyStatus_63_payload = debounce_1_keyStatus_63_payload;
  assign keyStatus_64_valid = debounce_1_keyStatus_64_valid;
  assign keyStatus_64_payload = debounce_1_keyStatus_64_payload;
  assign keyStatus_65_valid = debounce_1_keyStatus_65_valid;
  assign keyStatus_65_payload = debounce_1_keyStatus_65_payload;
  assign keyStatus_66_valid = debounce_1_keyStatus_66_valid;
  assign keyStatus_66_payload = debounce_1_keyStatus_66_payload;
  assign keyStatus_67_valid = debounce_1_keyStatus_67_valid;
  assign keyStatus_67_payload = debounce_1_keyStatus_67_payload;
  assign keyStatus_68_valid = debounce_1_keyStatus_68_valid;
  assign keyStatus_68_payload = debounce_1_keyStatus_68_payload;
  assign keyStatus_69_valid = debounce_1_keyStatus_69_valid;
  assign keyStatus_69_payload = debounce_1_keyStatus_69_payload;
  assign keyStatus_70_valid = debounce_1_keyStatus_70_valid;
  assign keyStatus_70_payload = debounce_1_keyStatus_70_payload;
  assign keyStatus_71_valid = debounce_1_keyStatus_71_valid;
  assign keyStatus_71_payload = debounce_1_keyStatus_71_payload;
  assign keyStatus_72_valid = debounce_1_keyStatus_72_valid;
  assign keyStatus_72_payload = debounce_1_keyStatus_72_payload;
  assign keyStatus_73_valid = debounce_1_keyStatus_73_valid;
  assign keyStatus_73_payload = debounce_1_keyStatus_73_payload;
  assign keyStatus_74_valid = debounce_1_keyStatus_74_valid;
  assign keyStatus_74_payload = debounce_1_keyStatus_74_payload;
  assign keyStatus_75_valid = debounce_1_keyStatus_75_valid;
  assign keyStatus_75_payload = debounce_1_keyStatus_75_payload;
  assign keyStatus_76_valid = debounce_1_keyStatus_76_valid;
  assign keyStatus_76_payload = debounce_1_keyStatus_76_payload;
  assign keyStatus_77_valid = debounce_1_keyStatus_77_valid;
  assign keyStatus_77_payload = debounce_1_keyStatus_77_payload;
  assign keyStatus_78_valid = debounce_1_keyStatus_78_valid;
  assign keyStatus_78_payload = debounce_1_keyStatus_78_payload;
  assign keyStatus_79_valid = debounce_1_keyStatus_79_valid;
  assign keyStatus_79_payload = debounce_1_keyStatus_79_payload;
  assign keyStatus_80_valid = debounce_1_keyStatus_80_valid;
  assign keyStatus_80_payload = debounce_1_keyStatus_80_payload;
  assign keyStatus_81_valid = debounce_1_keyStatus_81_valid;
  assign keyStatus_81_payload = debounce_1_keyStatus_81_payload;
  assign keyStatus_82_valid = debounce_1_keyStatus_82_valid;
  assign keyStatus_82_payload = debounce_1_keyStatus_82_payload;
  assign keyStatus_83_valid = debounce_1_keyStatus_83_valid;
  assign keyStatus_83_payload = debounce_1_keyStatus_83_payload;
  assign keyStatus_84_valid = debounce_1_keyStatus_84_valid;
  assign keyStatus_84_payload = debounce_1_keyStatus_84_payload;
  assign keyStatus_85_valid = debounce_1_keyStatus_85_valid;
  assign keyStatus_85_payload = debounce_1_keyStatus_85_payload;
  assign keyStatus_86_valid = debounce_1_keyStatus_86_valid;
  assign keyStatus_86_payload = debounce_1_keyStatus_86_payload;
  assign keyStatus_87_valid = debounce_1_keyStatus_87_valid;
  assign keyStatus_87_payload = debounce_1_keyStatus_87_payload;
  assign keyStatus_88_valid = debounce_1_keyStatus_88_valid;
  assign keyStatus_88_payload = debounce_1_keyStatus_88_payload;
  assign keyStatus_89_valid = debounce_1_keyStatus_89_valid;
  assign keyStatus_89_payload = debounce_1_keyStatus_89_payload;
  assign keyStatus_90_valid = debounce_1_keyStatus_90_valid;
  assign keyStatus_90_payload = debounce_1_keyStatus_90_payload;
  assign keyStatus_91_valid = debounce_1_keyStatus_91_valid;
  assign keyStatus_91_payload = debounce_1_keyStatus_91_payload;
  assign keyStatus_92_valid = debounce_1_keyStatus_92_valid;
  assign keyStatus_92_payload = debounce_1_keyStatus_92_payload;
  assign keyStatus_93_valid = debounce_1_keyStatus_93_valid;
  assign keyStatus_93_payload = debounce_1_keyStatus_93_payload;
  assign keyStatus_94_valid = debounce_1_keyStatus_94_valid;
  assign keyStatus_94_payload = debounce_1_keyStatus_94_payload;
  assign keyStatus_95_valid = debounce_1_keyStatus_95_valid;
  assign keyStatus_95_payload = debounce_1_keyStatus_95_payload;
  assign keyStatus_96_valid = debounce_1_keyStatus_96_valid;
  assign keyStatus_96_payload = debounce_1_keyStatus_96_payload;
  assign keyStatus_97_valid = debounce_1_keyStatus_97_valid;
  assign keyStatus_97_payload = debounce_1_keyStatus_97_payload;
  assign keyStatus_98_valid = debounce_1_keyStatus_98_valid;
  assign keyStatus_98_payload = debounce_1_keyStatus_98_payload;
  assign keyStatus_99_valid = debounce_1_keyStatus_99_valid;
  assign keyStatus_99_payload = debounce_1_keyStatus_99_payload;
  assign keyStatus_100_valid = debounce_1_keyStatus_100_valid;
  assign keyStatus_100_payload = debounce_1_keyStatus_100_payload;
  assign keyStatus_101_valid = debounce_1_keyStatus_101_valid;
  assign keyStatus_101_payload = debounce_1_keyStatus_101_payload;
  assign keyStatus_102_valid = debounce_1_keyStatus_102_valid;
  assign keyStatus_102_payload = debounce_1_keyStatus_102_payload;
  assign _zz_3 = (_zz_2 == 7'h60);
  assign _zz_7 = (_zz_6 == 7'h66);
  assign _zz_8 = (_zz_7 && _zz_4);
  always @ (*) begin
    if(_zz_8)begin
      _zz_5 = 7'h0;
    end else begin
      _zz_5 = (_zz_6 + _zz_14);
    end
    if(1'b0)begin
      _zz_5 = 7'h0;
    end
  end

  assign _zz_4 = 1'b1;
  assign scanIdx_valid = _zz_9;
  assign scanIdx_payload = {_zz_10,_zz_6};
  always @ (posedge CLK_50 or posedge _zz_1) begin
    if (_zz_1) begin
      clkScan_state <= 1'b0;
      clkScan_counter_value <= 11'h0;
      _zz_2 <= 7'h0;
      _zz_3_regNext <= 1'b0;
    end else begin
      clkScan_counter_value <= clkScan_counter_valueNext;
      if(clkScan_counter_willOverflow)begin
        clkScan_state <= 1'b1;
      end
      if(clkScan_state)begin
        clkScan_state <= 1'b0;
      end
      _zz_2 <= (_zz_2 + 7'h01);
      if(_zz_3)begin
        _zz_2 <= 7'h0;
      end
      _zz_3_regNext <= _zz_3;
    end
  end

  always @ (posedge CLK_50 or posedge _zz_1) begin
    if (_zz_1) begin
      _zz_6 <= 7'h0;
    end else begin
      if(_zz_3_regNext) begin
        _zz_6 <= _zz_5;
      end
    end
  end


endmodule

module BufferCC_1 (
  input               io_dataIn,
  output              io_dataOut,
  input               CLK_50,
  input               _zz_1
);
  (* async_reg = "true" *) reg                 buffers_0;
  (* async_reg = "true" *) reg                 buffers_1;

  assign io_dataOut = buffers_1;
  always @ (posedge CLK_50 or posedge _zz_1) begin
    if (_zz_1) begin
      buffers_0 <= 1'b1;
      buffers_1 <= 1'b1;
    end else begin
      buffers_0 <= io_dataIn;
      buffers_1 <= buffers_0;
    end
  end


endmodule

module ResetController (
  input               io_clock,
  input               io_externalReset,
  output              io_globalReset
);
  wire       [0:0]    _zz_14;
  wire       [15:0]   _zz_15;
  wire       [0:0]    _zz_16;
  wire       [27:0]   _zz_17;
  reg                 _zz_1;
  reg        [15:0]   _zz_2;
  reg        [15:0]   _zz_3 = 16'h0;
  wire                _zz_4;
  wire                _zz_5;
  reg                 _zz_6 = 1'b1;
  reg                 _zz_7;
  reg                 _zz_8;
  reg        [27:0]   _zz_9;
  reg        [27:0]   _zz_10 = 28'h0;
  wire                _zz_11;
  wire                _zz_12;
  reg                 io_externalReset_regNext = 1'b0;
  reg                 _zz_13;

  assign _zz_14 = _zz_1;
  assign _zz_15 = {15'd0, _zz_14};
  assign _zz_16 = _zz_7;
  assign _zz_17 = {27'd0, _zz_16};
  always @ (*) begin
    _zz_1 = 1'b0;
    if(_zz_6)begin
      _zz_1 = 1'b1;
    end
  end

  assign _zz_4 = (_zz_3 == 16'hc34f);
  assign _zz_5 = (_zz_4 && _zz_1);
  always @ (*) begin
    if(_zz_5)begin
      _zz_2 = 16'h0;
    end else begin
      _zz_2 = (_zz_3 + _zz_15);
    end
    if(1'b0)begin
      _zz_2 = 16'h0;
    end
  end

  always @ (*) begin
    _zz_7 = 1'b0;
    if(io_externalReset)begin
      _zz_7 = 1'b1;
    end
  end

  always @ (*) begin
    _zz_8 = 1'b0;
    if((io_externalReset && (! io_externalReset_regNext)))begin
      _zz_8 = 1'b1;
    end
  end

  assign _zz_11 = (_zz_10 == 28'h8f0d17f);
  assign _zz_12 = (_zz_11 && _zz_7);
  always @ (*) begin
    if(_zz_12)begin
      _zz_9 = 28'h0;
    end else begin
      _zz_9 = (_zz_10 + _zz_17);
    end
    if(_zz_8)begin
      _zz_9 = 28'h0;
    end
  end

  assign io_globalReset = _zz_13;
  always @ (posedge io_clock) begin
    _zz_3 <= _zz_2;
    if(_zz_4)begin
      _zz_6 <= 1'b0;
    end
    _zz_10 <= _zz_9;
    io_externalReset_regNext <= io_externalReset;
  end

  always @ (posedge io_clock) begin
    _zz_13 <= (_zz_6 || _zz_12);
  end


endmodule

module UartCtrl (
  input      [2:0]    io_config_frame_dataLength,
  input      `UartStopType_defaultEncoding_type io_config_frame_stop,
  input      `UartParityType_defaultEncoding_type io_config_frame_parity,
  input      [19:0]   io_config_clockDivider,
  input               io_write_valid,
  output reg          io_write_ready,
  input      [7:0]    io_write_payload,
  output              io_read_valid,
  input               io_read_ready,
  output     [7:0]    io_read_payload,
  output              io_uart_txd,
  input               io_uart_rxd,
  output              io_readError,
  input               io_writeBreak,
  output              io_readBreak,
  input               CLK_50,
  input               _zz_1
);
  wire                _zz_2;
  wire                tx_io_write_ready;
  wire                tx_io_txd;
  wire                rx_io_read_valid;
  wire       [7:0]    rx_io_read_payload;
  wire                rx_io_rts;
  wire                rx_io_error;
  wire                rx_io_break;
  reg        [19:0]   clockDivider_counter;
  wire                clockDivider_tick;
  reg                 io_write_thrown_valid;
  wire                io_write_thrown_ready;
  wire       [7:0]    io_write_thrown_payload;
  `ifndef SYNTHESIS
  reg [23:0] io_config_frame_stop_string;
  reg [31:0] io_config_frame_parity_string;
  `endif


  UartCtrlTx tx (
    .io_configFrame_dataLength    (io_config_frame_dataLength[2:0]  ), //i
    .io_configFrame_stop          (io_config_frame_stop             ), //i
    .io_configFrame_parity        (io_config_frame_parity[1:0]      ), //i
    .io_samplingTick              (clockDivider_tick                ), //i
    .io_write_valid               (io_write_thrown_valid            ), //i
    .io_write_ready               (tx_io_write_ready                ), //o
    .io_write_payload             (io_write_thrown_payload[7:0]     ), //i
    .io_cts                       (_zz_2                            ), //i
    .io_txd                       (tx_io_txd                        ), //o
    .io_break                     (io_writeBreak                    ), //i
    .CLK_50                       (CLK_50                           ), //i
    ._zz_2                        (_zz_1                            )  //i
  );
  UartCtrlRx rx (
    .io_configFrame_dataLength    (io_config_frame_dataLength[2:0]  ), //i
    .io_configFrame_stop          (io_config_frame_stop             ), //i
    .io_configFrame_parity        (io_config_frame_parity[1:0]      ), //i
    .io_samplingTick              (clockDivider_tick                ), //i
    .io_read_valid                (rx_io_read_valid                 ), //o
    .io_read_ready                (io_read_ready                    ), //i
    .io_read_payload              (rx_io_read_payload[7:0]          ), //o
    .io_rxd                       (io_uart_rxd                      ), //i
    .io_rts                       (rx_io_rts                        ), //o
    .io_error                     (rx_io_error                      ), //o
    .io_break                     (rx_io_break                      ), //o
    .CLK_50                       (CLK_50                           ), //i
    ._zz_2                        (_zz_1                            )  //i
  );
  `ifndef SYNTHESIS
  always @(*) begin
    case(io_config_frame_stop)
      `UartStopType_defaultEncoding_ONE : io_config_frame_stop_string = "ONE";
      `UartStopType_defaultEncoding_TWO : io_config_frame_stop_string = "TWO";
      default : io_config_frame_stop_string = "???";
    endcase
  end
  always @(*) begin
    case(io_config_frame_parity)
      `UartParityType_defaultEncoding_NONE : io_config_frame_parity_string = "NONE";
      `UartParityType_defaultEncoding_EVEN : io_config_frame_parity_string = "EVEN";
      `UartParityType_defaultEncoding_ODD : io_config_frame_parity_string = "ODD ";
      default : io_config_frame_parity_string = "????";
    endcase
  end
  `endif

  assign clockDivider_tick = (clockDivider_counter == 20'h0);
  always @ (*) begin
    io_write_thrown_valid = io_write_valid;
    if(rx_io_break)begin
      io_write_thrown_valid = 1'b0;
    end
  end

  always @ (*) begin
    io_write_ready = io_write_thrown_ready;
    if(rx_io_break)begin
      io_write_ready = 1'b1;
    end
  end

  assign io_write_thrown_payload = io_write_payload;
  assign io_write_thrown_ready = tx_io_write_ready;
  assign io_read_valid = rx_io_read_valid;
  assign io_read_payload = rx_io_read_payload;
  assign io_uart_txd = tx_io_txd;
  assign io_readError = rx_io_error;
  assign _zz_2 = 1'b0;
  assign io_readBreak = rx_io_break;
  always @ (posedge CLK_50 or posedge _zz_1) begin
    if (_zz_1) begin
      clockDivider_counter <= 20'h0;
    end else begin
      clockDivider_counter <= (clockDivider_counter - 20'h00001);
      if(clockDivider_tick)begin
        clockDivider_counter <= io_config_clockDivider;
      end
    end
  end


endmodule

module Debounce (
  input      [102:0]  key_down,
  output              keyStatus_0_valid,
  output              keyStatus_0_payload,
  output              keyStatus_1_valid,
  output              keyStatus_1_payload,
  output              keyStatus_2_valid,
  output              keyStatus_2_payload,
  output              keyStatus_3_valid,
  output              keyStatus_3_payload,
  output              keyStatus_4_valid,
  output              keyStatus_4_payload,
  output              keyStatus_5_valid,
  output              keyStatus_5_payload,
  output              keyStatus_6_valid,
  output              keyStatus_6_payload,
  output              keyStatus_7_valid,
  output              keyStatus_7_payload,
  output              keyStatus_8_valid,
  output              keyStatus_8_payload,
  output              keyStatus_9_valid,
  output              keyStatus_9_payload,
  output              keyStatus_10_valid,
  output              keyStatus_10_payload,
  output              keyStatus_11_valid,
  output              keyStatus_11_payload,
  output              keyStatus_12_valid,
  output              keyStatus_12_payload,
  output              keyStatus_13_valid,
  output              keyStatus_13_payload,
  output              keyStatus_14_valid,
  output              keyStatus_14_payload,
  output              keyStatus_15_valid,
  output              keyStatus_15_payload,
  output              keyStatus_16_valid,
  output              keyStatus_16_payload,
  output              keyStatus_17_valid,
  output              keyStatus_17_payload,
  output              keyStatus_18_valid,
  output              keyStatus_18_payload,
  output              keyStatus_19_valid,
  output              keyStatus_19_payload,
  output              keyStatus_20_valid,
  output              keyStatus_20_payload,
  output              keyStatus_21_valid,
  output              keyStatus_21_payload,
  output              keyStatus_22_valid,
  output              keyStatus_22_payload,
  output              keyStatus_23_valid,
  output              keyStatus_23_payload,
  output              keyStatus_24_valid,
  output              keyStatus_24_payload,
  output              keyStatus_25_valid,
  output              keyStatus_25_payload,
  output              keyStatus_26_valid,
  output              keyStatus_26_payload,
  output              keyStatus_27_valid,
  output              keyStatus_27_payload,
  output              keyStatus_28_valid,
  output              keyStatus_28_payload,
  output              keyStatus_29_valid,
  output              keyStatus_29_payload,
  output              keyStatus_30_valid,
  output              keyStatus_30_payload,
  output              keyStatus_31_valid,
  output              keyStatus_31_payload,
  output              keyStatus_32_valid,
  output              keyStatus_32_payload,
  output              keyStatus_33_valid,
  output              keyStatus_33_payload,
  output              keyStatus_34_valid,
  output              keyStatus_34_payload,
  output              keyStatus_35_valid,
  output              keyStatus_35_payload,
  output              keyStatus_36_valid,
  output              keyStatus_36_payload,
  output              keyStatus_37_valid,
  output              keyStatus_37_payload,
  output              keyStatus_38_valid,
  output              keyStatus_38_payload,
  output              keyStatus_39_valid,
  output              keyStatus_39_payload,
  output              keyStatus_40_valid,
  output              keyStatus_40_payload,
  output              keyStatus_41_valid,
  output              keyStatus_41_payload,
  output              keyStatus_42_valid,
  output              keyStatus_42_payload,
  output              keyStatus_43_valid,
  output              keyStatus_43_payload,
  output              keyStatus_44_valid,
  output              keyStatus_44_payload,
  output              keyStatus_45_valid,
  output              keyStatus_45_payload,
  output              keyStatus_46_valid,
  output              keyStatus_46_payload,
  output              keyStatus_47_valid,
  output              keyStatus_47_payload,
  output              keyStatus_48_valid,
  output              keyStatus_48_payload,
  output              keyStatus_49_valid,
  output              keyStatus_49_payload,
  output              keyStatus_50_valid,
  output              keyStatus_50_payload,
  output              keyStatus_51_valid,
  output              keyStatus_51_payload,
  output              keyStatus_52_valid,
  output              keyStatus_52_payload,
  output              keyStatus_53_valid,
  output              keyStatus_53_payload,
  output              keyStatus_54_valid,
  output              keyStatus_54_payload,
  output              keyStatus_55_valid,
  output              keyStatus_55_payload,
  output              keyStatus_56_valid,
  output              keyStatus_56_payload,
  output              keyStatus_57_valid,
  output              keyStatus_57_payload,
  output              keyStatus_58_valid,
  output              keyStatus_58_payload,
  output              keyStatus_59_valid,
  output              keyStatus_59_payload,
  output              keyStatus_60_valid,
  output              keyStatus_60_payload,
  output              keyStatus_61_valid,
  output              keyStatus_61_payload,
  output              keyStatus_62_valid,
  output              keyStatus_62_payload,
  output              keyStatus_63_valid,
  output              keyStatus_63_payload,
  output              keyStatus_64_valid,
  output              keyStatus_64_payload,
  output              keyStatus_65_valid,
  output              keyStatus_65_payload,
  output              keyStatus_66_valid,
  output              keyStatus_66_payload,
  output              keyStatus_67_valid,
  output              keyStatus_67_payload,
  output              keyStatus_68_valid,
  output              keyStatus_68_payload,
  output              keyStatus_69_valid,
  output              keyStatus_69_payload,
  output              keyStatus_70_valid,
  output              keyStatus_70_payload,
  output              keyStatus_71_valid,
  output              keyStatus_71_payload,
  output              keyStatus_72_valid,
  output              keyStatus_72_payload,
  output              keyStatus_73_valid,
  output              keyStatus_73_payload,
  output              keyStatus_74_valid,
  output              keyStatus_74_payload,
  output              keyStatus_75_valid,
  output              keyStatus_75_payload,
  output              keyStatus_76_valid,
  output              keyStatus_76_payload,
  output              keyStatus_77_valid,
  output              keyStatus_77_payload,
  output              keyStatus_78_valid,
  output              keyStatus_78_payload,
  output              keyStatus_79_valid,
  output              keyStatus_79_payload,
  output              keyStatus_80_valid,
  output              keyStatus_80_payload,
  output              keyStatus_81_valid,
  output              keyStatus_81_payload,
  output              keyStatus_82_valid,
  output              keyStatus_82_payload,
  output              keyStatus_83_valid,
  output              keyStatus_83_payload,
  output              keyStatus_84_valid,
  output              keyStatus_84_payload,
  output              keyStatus_85_valid,
  output              keyStatus_85_payload,
  output              keyStatus_86_valid,
  output              keyStatus_86_payload,
  output              keyStatus_87_valid,
  output              keyStatus_87_payload,
  output              keyStatus_88_valid,
  output              keyStatus_88_payload,
  output              keyStatus_89_valid,
  output              keyStatus_89_payload,
  output              keyStatus_90_valid,
  output              keyStatus_90_payload,
  output              keyStatus_91_valid,
  output              keyStatus_91_payload,
  output              keyStatus_92_valid,
  output              keyStatus_92_payload,
  output              keyStatus_93_valid,
  output              keyStatus_93_payload,
  output              keyStatus_94_valid,
  output              keyStatus_94_payload,
  output              keyStatus_95_valid,
  output              keyStatus_95_payload,
  output              keyStatus_96_valid,
  output              keyStatus_96_payload,
  output              keyStatus_97_valid,
  output              keyStatus_97_payload,
  output              keyStatus_98_valid,
  output              keyStatus_98_payload,
  output              keyStatus_99_valid,
  output              keyStatus_99_payload,
  output              keyStatus_100_valid,
  output              keyStatus_100_payload,
  output              keyStatus_101_valid,
  output              keyStatus_101_payload,
  output              keyStatus_102_valid,
  output              keyStatus_102_payload,
  input               CLK_50,
  input               _zz_3
);
  wire                _zz_4;
  wire                _zz_5;
  wire                _zz_6;
  wire                _zz_7;
  wire                _zz_8;
  wire                _zz_9;
  wire                _zz_10;
  wire                _zz_11;
  wire                _zz_12;
  wire                _zz_13;
  wire                _zz_14;
  wire                _zz_15;
  wire                _zz_16;
  wire                _zz_17;
  wire                _zz_18;
  wire                _zz_19;
  wire                _zz_20;
  wire                _zz_21;
  wire                _zz_22;
  wire                _zz_23;
  wire                _zz_24;
  wire                _zz_25;
  wire                _zz_26;
  wire                _zz_27;
  wire                _zz_28;
  wire                _zz_29;
  wire                _zz_30;
  wire                _zz_31;
  wire                _zz_32;
  wire                _zz_33;
  wire                _zz_34;
  wire                _zz_35;
  wire                _zz_36;
  wire                _zz_37;
  wire                _zz_38;
  wire                _zz_39;
  wire                _zz_40;
  wire                _zz_41;
  wire                _zz_42;
  wire                _zz_43;
  wire                _zz_44;
  wire                _zz_45;
  wire                _zz_46;
  wire                _zz_47;
  wire                _zz_48;
  wire                _zz_49;
  wire                _zz_50;
  wire                _zz_51;
  wire                _zz_52;
  wire                _zz_53;
  wire                _zz_54;
  wire                _zz_55;
  wire                _zz_56;
  wire                _zz_57;
  wire                _zz_58;
  wire                _zz_59;
  wire                _zz_60;
  wire                _zz_61;
  wire                _zz_62;
  wire                _zz_63;
  wire                _zz_64;
  wire                _zz_65;
  wire                _zz_66;
  wire                _zz_67;
  wire                _zz_68;
  wire                _zz_69;
  wire                _zz_70;
  wire                _zz_71;
  wire                _zz_72;
  wire                _zz_73;
  wire                _zz_74;
  wire                _zz_75;
  wire                _zz_76;
  wire                _zz_77;
  wire                _zz_78;
  wire                _zz_79;
  wire                _zz_80;
  wire                _zz_81;
  wire                _zz_82;
  wire                _zz_83;
  wire                _zz_84;
  wire                _zz_85;
  wire                _zz_86;
  wire                _zz_87;
  wire                _zz_88;
  wire                _zz_89;
  wire                _zz_90;
  wire                _zz_91;
  wire                _zz_92;
  wire                _zz_93;
  wire                _zz_94;
  wire                _zz_95;
  wire                _zz_96;
  wire                _zz_97;
  wire                _zz_98;
  wire                _zz_99;
  wire                _zz_100;
  wire                _zz_101;
  wire                _zz_102;
  wire                _zz_103;
  wire                _zz_104;
  wire                _zz_105;
  wire                _zz_106;
  wire                singleKey_103_filtered_valid;
  wire                singleKey_103_filtered_payload;
  wire                singleKey_104_filtered_valid;
  wire                singleKey_104_filtered_payload;
  wire                singleKey_105_filtered_valid;
  wire                singleKey_105_filtered_payload;
  wire                singleKey_106_filtered_valid;
  wire                singleKey_106_filtered_payload;
  wire                singleKey_107_filtered_valid;
  wire                singleKey_107_filtered_payload;
  wire                singleKey_108_filtered_valid;
  wire                singleKey_108_filtered_payload;
  wire                singleKey_109_filtered_valid;
  wire                singleKey_109_filtered_payload;
  wire                singleKey_110_filtered_valid;
  wire                singleKey_110_filtered_payload;
  wire                singleKey_111_filtered_valid;
  wire                singleKey_111_filtered_payload;
  wire                singleKey_112_filtered_valid;
  wire                singleKey_112_filtered_payload;
  wire                singleKey_113_filtered_valid;
  wire                singleKey_113_filtered_payload;
  wire                singleKey_114_filtered_valid;
  wire                singleKey_114_filtered_payload;
  wire                singleKey_115_filtered_valid;
  wire                singleKey_115_filtered_payload;
  wire                singleKey_116_filtered_valid;
  wire                singleKey_116_filtered_payload;
  wire                singleKey_117_filtered_valid;
  wire                singleKey_117_filtered_payload;
  wire                singleKey_118_filtered_valid;
  wire                singleKey_118_filtered_payload;
  wire                singleKey_119_filtered_valid;
  wire                singleKey_119_filtered_payload;
  wire                singleKey_120_filtered_valid;
  wire                singleKey_120_filtered_payload;
  wire                singleKey_121_filtered_valid;
  wire                singleKey_121_filtered_payload;
  wire                singleKey_122_filtered_valid;
  wire                singleKey_122_filtered_payload;
  wire                singleKey_123_filtered_valid;
  wire                singleKey_123_filtered_payload;
  wire                singleKey_124_filtered_valid;
  wire                singleKey_124_filtered_payload;
  wire                singleKey_125_filtered_valid;
  wire                singleKey_125_filtered_payload;
  wire                singleKey_126_filtered_valid;
  wire                singleKey_126_filtered_payload;
  wire                singleKey_127_filtered_valid;
  wire                singleKey_127_filtered_payload;
  wire                singleKey_128_filtered_valid;
  wire                singleKey_128_filtered_payload;
  wire                singleKey_129_filtered_valid;
  wire                singleKey_129_filtered_payload;
  wire                singleKey_130_filtered_valid;
  wire                singleKey_130_filtered_payload;
  wire                singleKey_131_filtered_valid;
  wire                singleKey_131_filtered_payload;
  wire                singleKey_132_filtered_valid;
  wire                singleKey_132_filtered_payload;
  wire                singleKey_133_filtered_valid;
  wire                singleKey_133_filtered_payload;
  wire                singleKey_134_filtered_valid;
  wire                singleKey_134_filtered_payload;
  wire                singleKey_135_filtered_valid;
  wire                singleKey_135_filtered_payload;
  wire                singleKey_136_filtered_valid;
  wire                singleKey_136_filtered_payload;
  wire                singleKey_137_filtered_valid;
  wire                singleKey_137_filtered_payload;
  wire                singleKey_138_filtered_valid;
  wire                singleKey_138_filtered_payload;
  wire                singleKey_139_filtered_valid;
  wire                singleKey_139_filtered_payload;
  wire                singleKey_140_filtered_valid;
  wire                singleKey_140_filtered_payload;
  wire                singleKey_141_filtered_valid;
  wire                singleKey_141_filtered_payload;
  wire                singleKey_142_filtered_valid;
  wire                singleKey_142_filtered_payload;
  wire                singleKey_143_filtered_valid;
  wire                singleKey_143_filtered_payload;
  wire                singleKey_144_filtered_valid;
  wire                singleKey_144_filtered_payload;
  wire                singleKey_145_filtered_valid;
  wire                singleKey_145_filtered_payload;
  wire                singleKey_146_filtered_valid;
  wire                singleKey_146_filtered_payload;
  wire                singleKey_147_filtered_valid;
  wire                singleKey_147_filtered_payload;
  wire                singleKey_148_filtered_valid;
  wire                singleKey_148_filtered_payload;
  wire                singleKey_149_filtered_valid;
  wire                singleKey_149_filtered_payload;
  wire                singleKey_150_filtered_valid;
  wire                singleKey_150_filtered_payload;
  wire                singleKey_151_filtered_valid;
  wire                singleKey_151_filtered_payload;
  wire                singleKey_152_filtered_valid;
  wire                singleKey_152_filtered_payload;
  wire                singleKey_153_filtered_valid;
  wire                singleKey_153_filtered_payload;
  wire                singleKey_154_filtered_valid;
  wire                singleKey_154_filtered_payload;
  wire                singleKey_155_filtered_valid;
  wire                singleKey_155_filtered_payload;
  wire                singleKey_156_filtered_valid;
  wire                singleKey_156_filtered_payload;
  wire                singleKey_157_filtered_valid;
  wire                singleKey_157_filtered_payload;
  wire                singleKey_158_filtered_valid;
  wire                singleKey_158_filtered_payload;
  wire                singleKey_159_filtered_valid;
  wire                singleKey_159_filtered_payload;
  wire                singleKey_160_filtered_valid;
  wire                singleKey_160_filtered_payload;
  wire                singleKey_161_filtered_valid;
  wire                singleKey_161_filtered_payload;
  wire                singleKey_162_filtered_valid;
  wire                singleKey_162_filtered_payload;
  wire                singleKey_163_filtered_valid;
  wire                singleKey_163_filtered_payload;
  wire                singleKey_164_filtered_valid;
  wire                singleKey_164_filtered_payload;
  wire                singleKey_165_filtered_valid;
  wire                singleKey_165_filtered_payload;
  wire                singleKey_166_filtered_valid;
  wire                singleKey_166_filtered_payload;
  wire                singleKey_167_filtered_valid;
  wire                singleKey_167_filtered_payload;
  wire                singleKey_168_filtered_valid;
  wire                singleKey_168_filtered_payload;
  wire                singleKey_169_filtered_valid;
  wire                singleKey_169_filtered_payload;
  wire                singleKey_170_filtered_valid;
  wire                singleKey_170_filtered_payload;
  wire                singleKey_171_filtered_valid;
  wire                singleKey_171_filtered_payload;
  wire                singleKey_172_filtered_valid;
  wire                singleKey_172_filtered_payload;
  wire                singleKey_173_filtered_valid;
  wire                singleKey_173_filtered_payload;
  wire                singleKey_174_filtered_valid;
  wire                singleKey_174_filtered_payload;
  wire                singleKey_175_filtered_valid;
  wire                singleKey_175_filtered_payload;
  wire                singleKey_176_filtered_valid;
  wire                singleKey_176_filtered_payload;
  wire                singleKey_177_filtered_valid;
  wire                singleKey_177_filtered_payload;
  wire                singleKey_178_filtered_valid;
  wire                singleKey_178_filtered_payload;
  wire                singleKey_179_filtered_valid;
  wire                singleKey_179_filtered_payload;
  wire                singleKey_180_filtered_valid;
  wire                singleKey_180_filtered_payload;
  wire                singleKey_181_filtered_valid;
  wire                singleKey_181_filtered_payload;
  wire                singleKey_182_filtered_valid;
  wire                singleKey_182_filtered_payload;
  wire                singleKey_183_filtered_valid;
  wire                singleKey_183_filtered_payload;
  wire                singleKey_184_filtered_valid;
  wire                singleKey_184_filtered_payload;
  wire                singleKey_185_filtered_valid;
  wire                singleKey_185_filtered_payload;
  wire                singleKey_186_filtered_valid;
  wire                singleKey_186_filtered_payload;
  wire                singleKey_187_filtered_valid;
  wire                singleKey_187_filtered_payload;
  wire                singleKey_188_filtered_valid;
  wire                singleKey_188_filtered_payload;
  wire                singleKey_189_filtered_valid;
  wire                singleKey_189_filtered_payload;
  wire                singleKey_190_filtered_valid;
  wire                singleKey_190_filtered_payload;
  wire                singleKey_191_filtered_valid;
  wire                singleKey_191_filtered_payload;
  wire                singleKey_192_filtered_valid;
  wire                singleKey_192_filtered_payload;
  wire                singleKey_193_filtered_valid;
  wire                singleKey_193_filtered_payload;
  wire                singleKey_194_filtered_valid;
  wire                singleKey_194_filtered_payload;
  wire                singleKey_195_filtered_valid;
  wire                singleKey_195_filtered_payload;
  wire                singleKey_196_filtered_valid;
  wire                singleKey_196_filtered_payload;
  wire                singleKey_197_filtered_valid;
  wire                singleKey_197_filtered_payload;
  wire                singleKey_198_filtered_valid;
  wire                singleKey_198_filtered_payload;
  wire                singleKey_199_filtered_valid;
  wire                singleKey_199_filtered_payload;
  wire                singleKey_200_filtered_valid;
  wire                singleKey_200_filtered_payload;
  wire                singleKey_201_filtered_valid;
  wire                singleKey_201_filtered_payload;
  wire                singleKey_202_filtered_valid;
  wire                singleKey_202_filtered_payload;
  wire                singleKey_203_filtered_valid;
  wire                singleKey_203_filtered_payload;
  wire                singleKey_204_filtered_valid;
  wire                singleKey_204_filtered_payload;
  wire                singleKey_205_filtered_valid;
  wire                singleKey_205_filtered_payload;
  reg        [13:0]   _zz_1;
  wire                _zz_2;
  reg                 _zz_2_regNext;

  SingleKey singleKey_103 (
    .raw                 (_zz_4                           ), //i
    .filtered_valid      (singleKey_103_filtered_valid    ), //o
    .filtered_payload    (singleKey_103_filtered_payload  ), //o
    .CLK_50              (CLK_50                          ), //i
    ._zz_3               (_zz_3                           ), //i
    ._zz_4               (_zz_2_regNext                   )  //i
  );
  SingleKey singleKey_104 (
    .raw                 (_zz_5                           ), //i
    .filtered_valid      (singleKey_104_filtered_valid    ), //o
    .filtered_payload    (singleKey_104_filtered_payload  ), //o
    .CLK_50              (CLK_50                          ), //i
    ._zz_3               (_zz_3                           ), //i
    ._zz_4               (_zz_2_regNext                   )  //i
  );
  SingleKey singleKey_105 (
    .raw                 (_zz_6                           ), //i
    .filtered_valid      (singleKey_105_filtered_valid    ), //o
    .filtered_payload    (singleKey_105_filtered_payload  ), //o
    .CLK_50              (CLK_50                          ), //i
    ._zz_3               (_zz_3                           ), //i
    ._zz_4               (_zz_2_regNext                   )  //i
  );
  SingleKey singleKey_106 (
    .raw                 (_zz_7                           ), //i
    .filtered_valid      (singleKey_106_filtered_valid    ), //o
    .filtered_payload    (singleKey_106_filtered_payload  ), //o
    .CLK_50              (CLK_50                          ), //i
    ._zz_3               (_zz_3                           ), //i
    ._zz_4               (_zz_2_regNext                   )  //i
  );
  SingleKey singleKey_107 (
    .raw                 (_zz_8                           ), //i
    .filtered_valid      (singleKey_107_filtered_valid    ), //o
    .filtered_payload    (singleKey_107_filtered_payload  ), //o
    .CLK_50              (CLK_50                          ), //i
    ._zz_3               (_zz_3                           ), //i
    ._zz_4               (_zz_2_regNext                   )  //i
  );
  SingleKey singleKey_108 (
    .raw                 (_zz_9                           ), //i
    .filtered_valid      (singleKey_108_filtered_valid    ), //o
    .filtered_payload    (singleKey_108_filtered_payload  ), //o
    .CLK_50              (CLK_50                          ), //i
    ._zz_3               (_zz_3                           ), //i
    ._zz_4               (_zz_2_regNext                   )  //i
  );
  SingleKey singleKey_109 (
    .raw                 (_zz_10                          ), //i
    .filtered_valid      (singleKey_109_filtered_valid    ), //o
    .filtered_payload    (singleKey_109_filtered_payload  ), //o
    .CLK_50              (CLK_50                          ), //i
    ._zz_3               (_zz_3                           ), //i
    ._zz_4               (_zz_2_regNext                   )  //i
  );
  SingleKey singleKey_110 (
    .raw                 (_zz_11                          ), //i
    .filtered_valid      (singleKey_110_filtered_valid    ), //o
    .filtered_payload    (singleKey_110_filtered_payload  ), //o
    .CLK_50              (CLK_50                          ), //i
    ._zz_3               (_zz_3                           ), //i
    ._zz_4               (_zz_2_regNext                   )  //i
  );
  SingleKey singleKey_111 (
    .raw                 (_zz_12                          ), //i
    .filtered_valid      (singleKey_111_filtered_valid    ), //o
    .filtered_payload    (singleKey_111_filtered_payload  ), //o
    .CLK_50              (CLK_50                          ), //i
    ._zz_3               (_zz_3                           ), //i
    ._zz_4               (_zz_2_regNext                   )  //i
  );
  SingleKey singleKey_112 (
    .raw                 (_zz_13                          ), //i
    .filtered_valid      (singleKey_112_filtered_valid    ), //o
    .filtered_payload    (singleKey_112_filtered_payload  ), //o
    .CLK_50              (CLK_50                          ), //i
    ._zz_3               (_zz_3                           ), //i
    ._zz_4               (_zz_2_regNext                   )  //i
  );
  SingleKey singleKey_113 (
    .raw                 (_zz_14                          ), //i
    .filtered_valid      (singleKey_113_filtered_valid    ), //o
    .filtered_payload    (singleKey_113_filtered_payload  ), //o
    .CLK_50              (CLK_50                          ), //i
    ._zz_3               (_zz_3                           ), //i
    ._zz_4               (_zz_2_regNext                   )  //i
  );
  SingleKey singleKey_114 (
    .raw                 (_zz_15                          ), //i
    .filtered_valid      (singleKey_114_filtered_valid    ), //o
    .filtered_payload    (singleKey_114_filtered_payload  ), //o
    .CLK_50              (CLK_50                          ), //i
    ._zz_3               (_zz_3                           ), //i
    ._zz_4               (_zz_2_regNext                   )  //i
  );
  SingleKey singleKey_115 (
    .raw                 (_zz_16                          ), //i
    .filtered_valid      (singleKey_115_filtered_valid    ), //o
    .filtered_payload    (singleKey_115_filtered_payload  ), //o
    .CLK_50              (CLK_50                          ), //i
    ._zz_3               (_zz_3                           ), //i
    ._zz_4               (_zz_2_regNext                   )  //i
  );
  SingleKey singleKey_116 (
    .raw                 (_zz_17                          ), //i
    .filtered_valid      (singleKey_116_filtered_valid    ), //o
    .filtered_payload    (singleKey_116_filtered_payload  ), //o
    .CLK_50              (CLK_50                          ), //i
    ._zz_3               (_zz_3                           ), //i
    ._zz_4               (_zz_2_regNext                   )  //i
  );
  SingleKey singleKey_117 (
    .raw                 (_zz_18                          ), //i
    .filtered_valid      (singleKey_117_filtered_valid    ), //o
    .filtered_payload    (singleKey_117_filtered_payload  ), //o
    .CLK_50              (CLK_50                          ), //i
    ._zz_3               (_zz_3                           ), //i
    ._zz_4               (_zz_2_regNext                   )  //i
  );
  SingleKey singleKey_118 (
    .raw                 (_zz_19                          ), //i
    .filtered_valid      (singleKey_118_filtered_valid    ), //o
    .filtered_payload    (singleKey_118_filtered_payload  ), //o
    .CLK_50              (CLK_50                          ), //i
    ._zz_3               (_zz_3                           ), //i
    ._zz_4               (_zz_2_regNext                   )  //i
  );
  SingleKey singleKey_119 (
    .raw                 (_zz_20                          ), //i
    .filtered_valid      (singleKey_119_filtered_valid    ), //o
    .filtered_payload    (singleKey_119_filtered_payload  ), //o
    .CLK_50              (CLK_50                          ), //i
    ._zz_3               (_zz_3                           ), //i
    ._zz_4               (_zz_2_regNext                   )  //i
  );
  SingleKey singleKey_120 (
    .raw                 (_zz_21                          ), //i
    .filtered_valid      (singleKey_120_filtered_valid    ), //o
    .filtered_payload    (singleKey_120_filtered_payload  ), //o
    .CLK_50              (CLK_50                          ), //i
    ._zz_3               (_zz_3                           ), //i
    ._zz_4               (_zz_2_regNext                   )  //i
  );
  SingleKey singleKey_121 (
    .raw                 (_zz_22                          ), //i
    .filtered_valid      (singleKey_121_filtered_valid    ), //o
    .filtered_payload    (singleKey_121_filtered_payload  ), //o
    .CLK_50              (CLK_50                          ), //i
    ._zz_3               (_zz_3                           ), //i
    ._zz_4               (_zz_2_regNext                   )  //i
  );
  SingleKey singleKey_122 (
    .raw                 (_zz_23                          ), //i
    .filtered_valid      (singleKey_122_filtered_valid    ), //o
    .filtered_payload    (singleKey_122_filtered_payload  ), //o
    .CLK_50              (CLK_50                          ), //i
    ._zz_3               (_zz_3                           ), //i
    ._zz_4               (_zz_2_regNext                   )  //i
  );
  SingleKey singleKey_123 (
    .raw                 (_zz_24                          ), //i
    .filtered_valid      (singleKey_123_filtered_valid    ), //o
    .filtered_payload    (singleKey_123_filtered_payload  ), //o
    .CLK_50              (CLK_50                          ), //i
    ._zz_3               (_zz_3                           ), //i
    ._zz_4               (_zz_2_regNext                   )  //i
  );
  SingleKey singleKey_124 (
    .raw                 (_zz_25                          ), //i
    .filtered_valid      (singleKey_124_filtered_valid    ), //o
    .filtered_payload    (singleKey_124_filtered_payload  ), //o
    .CLK_50              (CLK_50                          ), //i
    ._zz_3               (_zz_3                           ), //i
    ._zz_4               (_zz_2_regNext                   )  //i
  );
  SingleKey singleKey_125 (
    .raw                 (_zz_26                          ), //i
    .filtered_valid      (singleKey_125_filtered_valid    ), //o
    .filtered_payload    (singleKey_125_filtered_payload  ), //o
    .CLK_50              (CLK_50                          ), //i
    ._zz_3               (_zz_3                           ), //i
    ._zz_4               (_zz_2_regNext                   )  //i
  );
  SingleKey singleKey_126 (
    .raw                 (_zz_27                          ), //i
    .filtered_valid      (singleKey_126_filtered_valid    ), //o
    .filtered_payload    (singleKey_126_filtered_payload  ), //o
    .CLK_50              (CLK_50                          ), //i
    ._zz_3               (_zz_3                           ), //i
    ._zz_4               (_zz_2_regNext                   )  //i
  );
  SingleKey singleKey_127 (
    .raw                 (_zz_28                          ), //i
    .filtered_valid      (singleKey_127_filtered_valid    ), //o
    .filtered_payload    (singleKey_127_filtered_payload  ), //o
    .CLK_50              (CLK_50                          ), //i
    ._zz_3               (_zz_3                           ), //i
    ._zz_4               (_zz_2_regNext                   )  //i
  );
  SingleKey singleKey_128 (
    .raw                 (_zz_29                          ), //i
    .filtered_valid      (singleKey_128_filtered_valid    ), //o
    .filtered_payload    (singleKey_128_filtered_payload  ), //o
    .CLK_50              (CLK_50                          ), //i
    ._zz_3               (_zz_3                           ), //i
    ._zz_4               (_zz_2_regNext                   )  //i
  );
  SingleKey singleKey_129 (
    .raw                 (_zz_30                          ), //i
    .filtered_valid      (singleKey_129_filtered_valid    ), //o
    .filtered_payload    (singleKey_129_filtered_payload  ), //o
    .CLK_50              (CLK_50                          ), //i
    ._zz_3               (_zz_3                           ), //i
    ._zz_4               (_zz_2_regNext                   )  //i
  );
  SingleKey singleKey_130 (
    .raw                 (_zz_31                          ), //i
    .filtered_valid      (singleKey_130_filtered_valid    ), //o
    .filtered_payload    (singleKey_130_filtered_payload  ), //o
    .CLK_50              (CLK_50                          ), //i
    ._zz_3               (_zz_3                           ), //i
    ._zz_4               (_zz_2_regNext                   )  //i
  );
  SingleKey singleKey_131 (
    .raw                 (_zz_32                          ), //i
    .filtered_valid      (singleKey_131_filtered_valid    ), //o
    .filtered_payload    (singleKey_131_filtered_payload  ), //o
    .CLK_50              (CLK_50                          ), //i
    ._zz_3               (_zz_3                           ), //i
    ._zz_4               (_zz_2_regNext                   )  //i
  );
  SingleKey singleKey_132 (
    .raw                 (_zz_33                          ), //i
    .filtered_valid      (singleKey_132_filtered_valid    ), //o
    .filtered_payload    (singleKey_132_filtered_payload  ), //o
    .CLK_50              (CLK_50                          ), //i
    ._zz_3               (_zz_3                           ), //i
    ._zz_4               (_zz_2_regNext                   )  //i
  );
  SingleKey singleKey_133 (
    .raw                 (_zz_34                          ), //i
    .filtered_valid      (singleKey_133_filtered_valid    ), //o
    .filtered_payload    (singleKey_133_filtered_payload  ), //o
    .CLK_50              (CLK_50                          ), //i
    ._zz_3               (_zz_3                           ), //i
    ._zz_4               (_zz_2_regNext                   )  //i
  );
  SingleKey singleKey_134 (
    .raw                 (_zz_35                          ), //i
    .filtered_valid      (singleKey_134_filtered_valid    ), //o
    .filtered_payload    (singleKey_134_filtered_payload  ), //o
    .CLK_50              (CLK_50                          ), //i
    ._zz_3               (_zz_3                           ), //i
    ._zz_4               (_zz_2_regNext                   )  //i
  );
  SingleKey singleKey_135 (
    .raw                 (_zz_36                          ), //i
    .filtered_valid      (singleKey_135_filtered_valid    ), //o
    .filtered_payload    (singleKey_135_filtered_payload  ), //o
    .CLK_50              (CLK_50                          ), //i
    ._zz_3               (_zz_3                           ), //i
    ._zz_4               (_zz_2_regNext                   )  //i
  );
  SingleKey singleKey_136 (
    .raw                 (_zz_37                          ), //i
    .filtered_valid      (singleKey_136_filtered_valid    ), //o
    .filtered_payload    (singleKey_136_filtered_payload  ), //o
    .CLK_50              (CLK_50                          ), //i
    ._zz_3               (_zz_3                           ), //i
    ._zz_4               (_zz_2_regNext                   )  //i
  );
  SingleKey singleKey_137 (
    .raw                 (_zz_38                          ), //i
    .filtered_valid      (singleKey_137_filtered_valid    ), //o
    .filtered_payload    (singleKey_137_filtered_payload  ), //o
    .CLK_50              (CLK_50                          ), //i
    ._zz_3               (_zz_3                           ), //i
    ._zz_4               (_zz_2_regNext                   )  //i
  );
  SingleKey singleKey_138 (
    .raw                 (_zz_39                          ), //i
    .filtered_valid      (singleKey_138_filtered_valid    ), //o
    .filtered_payload    (singleKey_138_filtered_payload  ), //o
    .CLK_50              (CLK_50                          ), //i
    ._zz_3               (_zz_3                           ), //i
    ._zz_4               (_zz_2_regNext                   )  //i
  );
  SingleKey singleKey_139 (
    .raw                 (_zz_40                          ), //i
    .filtered_valid      (singleKey_139_filtered_valid    ), //o
    .filtered_payload    (singleKey_139_filtered_payload  ), //o
    .CLK_50              (CLK_50                          ), //i
    ._zz_3               (_zz_3                           ), //i
    ._zz_4               (_zz_2_regNext                   )  //i
  );
  SingleKey singleKey_140 (
    .raw                 (_zz_41                          ), //i
    .filtered_valid      (singleKey_140_filtered_valid    ), //o
    .filtered_payload    (singleKey_140_filtered_payload  ), //o
    .CLK_50              (CLK_50                          ), //i
    ._zz_3               (_zz_3                           ), //i
    ._zz_4               (_zz_2_regNext                   )  //i
  );
  SingleKey singleKey_141 (
    .raw                 (_zz_42                          ), //i
    .filtered_valid      (singleKey_141_filtered_valid    ), //o
    .filtered_payload    (singleKey_141_filtered_payload  ), //o
    .CLK_50              (CLK_50                          ), //i
    ._zz_3               (_zz_3                           ), //i
    ._zz_4               (_zz_2_regNext                   )  //i
  );
  SingleKey singleKey_142 (
    .raw                 (_zz_43                          ), //i
    .filtered_valid      (singleKey_142_filtered_valid    ), //o
    .filtered_payload    (singleKey_142_filtered_payload  ), //o
    .CLK_50              (CLK_50                          ), //i
    ._zz_3               (_zz_3                           ), //i
    ._zz_4               (_zz_2_regNext                   )  //i
  );
  SingleKey singleKey_143 (
    .raw                 (_zz_44                          ), //i
    .filtered_valid      (singleKey_143_filtered_valid    ), //o
    .filtered_payload    (singleKey_143_filtered_payload  ), //o
    .CLK_50              (CLK_50                          ), //i
    ._zz_3               (_zz_3                           ), //i
    ._zz_4               (_zz_2_regNext                   )  //i
  );
  SingleKey singleKey_144 (
    .raw                 (_zz_45                          ), //i
    .filtered_valid      (singleKey_144_filtered_valid    ), //o
    .filtered_payload    (singleKey_144_filtered_payload  ), //o
    .CLK_50              (CLK_50                          ), //i
    ._zz_3               (_zz_3                           ), //i
    ._zz_4               (_zz_2_regNext                   )  //i
  );
  SingleKey singleKey_145 (
    .raw                 (_zz_46                          ), //i
    .filtered_valid      (singleKey_145_filtered_valid    ), //o
    .filtered_payload    (singleKey_145_filtered_payload  ), //o
    .CLK_50              (CLK_50                          ), //i
    ._zz_3               (_zz_3                           ), //i
    ._zz_4               (_zz_2_regNext                   )  //i
  );
  SingleKey singleKey_146 (
    .raw                 (_zz_47                          ), //i
    .filtered_valid      (singleKey_146_filtered_valid    ), //o
    .filtered_payload    (singleKey_146_filtered_payload  ), //o
    .CLK_50              (CLK_50                          ), //i
    ._zz_3               (_zz_3                           ), //i
    ._zz_4               (_zz_2_regNext                   )  //i
  );
  SingleKey singleKey_147 (
    .raw                 (_zz_48                          ), //i
    .filtered_valid      (singleKey_147_filtered_valid    ), //o
    .filtered_payload    (singleKey_147_filtered_payload  ), //o
    .CLK_50              (CLK_50                          ), //i
    ._zz_3               (_zz_3                           ), //i
    ._zz_4               (_zz_2_regNext                   )  //i
  );
  SingleKey singleKey_148 (
    .raw                 (_zz_49                          ), //i
    .filtered_valid      (singleKey_148_filtered_valid    ), //o
    .filtered_payload    (singleKey_148_filtered_payload  ), //o
    .CLK_50              (CLK_50                          ), //i
    ._zz_3               (_zz_3                           ), //i
    ._zz_4               (_zz_2_regNext                   )  //i
  );
  SingleKey singleKey_149 (
    .raw                 (_zz_50                          ), //i
    .filtered_valid      (singleKey_149_filtered_valid    ), //o
    .filtered_payload    (singleKey_149_filtered_payload  ), //o
    .CLK_50              (CLK_50                          ), //i
    ._zz_3               (_zz_3                           ), //i
    ._zz_4               (_zz_2_regNext                   )  //i
  );
  SingleKey singleKey_150 (
    .raw                 (_zz_51                          ), //i
    .filtered_valid      (singleKey_150_filtered_valid    ), //o
    .filtered_payload    (singleKey_150_filtered_payload  ), //o
    .CLK_50              (CLK_50                          ), //i
    ._zz_3               (_zz_3                           ), //i
    ._zz_4               (_zz_2_regNext                   )  //i
  );
  SingleKey singleKey_151 (
    .raw                 (_zz_52                          ), //i
    .filtered_valid      (singleKey_151_filtered_valid    ), //o
    .filtered_payload    (singleKey_151_filtered_payload  ), //o
    .CLK_50              (CLK_50                          ), //i
    ._zz_3               (_zz_3                           ), //i
    ._zz_4               (_zz_2_regNext                   )  //i
  );
  SingleKey singleKey_152 (
    .raw                 (_zz_53                          ), //i
    .filtered_valid      (singleKey_152_filtered_valid    ), //o
    .filtered_payload    (singleKey_152_filtered_payload  ), //o
    .CLK_50              (CLK_50                          ), //i
    ._zz_3               (_zz_3                           ), //i
    ._zz_4               (_zz_2_regNext                   )  //i
  );
  SingleKey singleKey_153 (
    .raw                 (_zz_54                          ), //i
    .filtered_valid      (singleKey_153_filtered_valid    ), //o
    .filtered_payload    (singleKey_153_filtered_payload  ), //o
    .CLK_50              (CLK_50                          ), //i
    ._zz_3               (_zz_3                           ), //i
    ._zz_4               (_zz_2_regNext                   )  //i
  );
  SingleKey singleKey_154 (
    .raw                 (_zz_55                          ), //i
    .filtered_valid      (singleKey_154_filtered_valid    ), //o
    .filtered_payload    (singleKey_154_filtered_payload  ), //o
    .CLK_50              (CLK_50                          ), //i
    ._zz_3               (_zz_3                           ), //i
    ._zz_4               (_zz_2_regNext                   )  //i
  );
  SingleKey singleKey_155 (
    .raw                 (_zz_56                          ), //i
    .filtered_valid      (singleKey_155_filtered_valid    ), //o
    .filtered_payload    (singleKey_155_filtered_payload  ), //o
    .CLK_50              (CLK_50                          ), //i
    ._zz_3               (_zz_3                           ), //i
    ._zz_4               (_zz_2_regNext                   )  //i
  );
  SingleKey singleKey_156 (
    .raw                 (_zz_57                          ), //i
    .filtered_valid      (singleKey_156_filtered_valid    ), //o
    .filtered_payload    (singleKey_156_filtered_payload  ), //o
    .CLK_50              (CLK_50                          ), //i
    ._zz_3               (_zz_3                           ), //i
    ._zz_4               (_zz_2_regNext                   )  //i
  );
  SingleKey singleKey_157 (
    .raw                 (_zz_58                          ), //i
    .filtered_valid      (singleKey_157_filtered_valid    ), //o
    .filtered_payload    (singleKey_157_filtered_payload  ), //o
    .CLK_50              (CLK_50                          ), //i
    ._zz_3               (_zz_3                           ), //i
    ._zz_4               (_zz_2_regNext                   )  //i
  );
  SingleKey singleKey_158 (
    .raw                 (_zz_59                          ), //i
    .filtered_valid      (singleKey_158_filtered_valid    ), //o
    .filtered_payload    (singleKey_158_filtered_payload  ), //o
    .CLK_50              (CLK_50                          ), //i
    ._zz_3               (_zz_3                           ), //i
    ._zz_4               (_zz_2_regNext                   )  //i
  );
  SingleKey singleKey_159 (
    .raw                 (_zz_60                          ), //i
    .filtered_valid      (singleKey_159_filtered_valid    ), //o
    .filtered_payload    (singleKey_159_filtered_payload  ), //o
    .CLK_50              (CLK_50                          ), //i
    ._zz_3               (_zz_3                           ), //i
    ._zz_4               (_zz_2_regNext                   )  //i
  );
  SingleKey singleKey_160 (
    .raw                 (_zz_61                          ), //i
    .filtered_valid      (singleKey_160_filtered_valid    ), //o
    .filtered_payload    (singleKey_160_filtered_payload  ), //o
    .CLK_50              (CLK_50                          ), //i
    ._zz_3               (_zz_3                           ), //i
    ._zz_4               (_zz_2_regNext                   )  //i
  );
  SingleKey singleKey_161 (
    .raw                 (_zz_62                          ), //i
    .filtered_valid      (singleKey_161_filtered_valid    ), //o
    .filtered_payload    (singleKey_161_filtered_payload  ), //o
    .CLK_50              (CLK_50                          ), //i
    ._zz_3               (_zz_3                           ), //i
    ._zz_4               (_zz_2_regNext                   )  //i
  );
  SingleKey singleKey_162 (
    .raw                 (_zz_63                          ), //i
    .filtered_valid      (singleKey_162_filtered_valid    ), //o
    .filtered_payload    (singleKey_162_filtered_payload  ), //o
    .CLK_50              (CLK_50                          ), //i
    ._zz_3               (_zz_3                           ), //i
    ._zz_4               (_zz_2_regNext                   )  //i
  );
  SingleKey singleKey_163 (
    .raw                 (_zz_64                          ), //i
    .filtered_valid      (singleKey_163_filtered_valid    ), //o
    .filtered_payload    (singleKey_163_filtered_payload  ), //o
    .CLK_50              (CLK_50                          ), //i
    ._zz_3               (_zz_3                           ), //i
    ._zz_4               (_zz_2_regNext                   )  //i
  );
  SingleKey singleKey_164 (
    .raw                 (_zz_65                          ), //i
    .filtered_valid      (singleKey_164_filtered_valid    ), //o
    .filtered_payload    (singleKey_164_filtered_payload  ), //o
    .CLK_50              (CLK_50                          ), //i
    ._zz_3               (_zz_3                           ), //i
    ._zz_4               (_zz_2_regNext                   )  //i
  );
  SingleKey singleKey_165 (
    .raw                 (_zz_66                          ), //i
    .filtered_valid      (singleKey_165_filtered_valid    ), //o
    .filtered_payload    (singleKey_165_filtered_payload  ), //o
    .CLK_50              (CLK_50                          ), //i
    ._zz_3               (_zz_3                           ), //i
    ._zz_4               (_zz_2_regNext                   )  //i
  );
  SingleKey singleKey_166 (
    .raw                 (_zz_67                          ), //i
    .filtered_valid      (singleKey_166_filtered_valid    ), //o
    .filtered_payload    (singleKey_166_filtered_payload  ), //o
    .CLK_50              (CLK_50                          ), //i
    ._zz_3               (_zz_3                           ), //i
    ._zz_4               (_zz_2_regNext                   )  //i
  );
  SingleKey singleKey_167 (
    .raw                 (_zz_68                          ), //i
    .filtered_valid      (singleKey_167_filtered_valid    ), //o
    .filtered_payload    (singleKey_167_filtered_payload  ), //o
    .CLK_50              (CLK_50                          ), //i
    ._zz_3               (_zz_3                           ), //i
    ._zz_4               (_zz_2_regNext                   )  //i
  );
  SingleKey singleKey_168 (
    .raw                 (_zz_69                          ), //i
    .filtered_valid      (singleKey_168_filtered_valid    ), //o
    .filtered_payload    (singleKey_168_filtered_payload  ), //o
    .CLK_50              (CLK_50                          ), //i
    ._zz_3               (_zz_3                           ), //i
    ._zz_4               (_zz_2_regNext                   )  //i
  );
  SingleKey singleKey_169 (
    .raw                 (_zz_70                          ), //i
    .filtered_valid      (singleKey_169_filtered_valid    ), //o
    .filtered_payload    (singleKey_169_filtered_payload  ), //o
    .CLK_50              (CLK_50                          ), //i
    ._zz_3               (_zz_3                           ), //i
    ._zz_4               (_zz_2_regNext                   )  //i
  );
  SingleKey singleKey_170 (
    .raw                 (_zz_71                          ), //i
    .filtered_valid      (singleKey_170_filtered_valid    ), //o
    .filtered_payload    (singleKey_170_filtered_payload  ), //o
    .CLK_50              (CLK_50                          ), //i
    ._zz_3               (_zz_3                           ), //i
    ._zz_4               (_zz_2_regNext                   )  //i
  );
  SingleKey singleKey_171 (
    .raw                 (_zz_72                          ), //i
    .filtered_valid      (singleKey_171_filtered_valid    ), //o
    .filtered_payload    (singleKey_171_filtered_payload  ), //o
    .CLK_50              (CLK_50                          ), //i
    ._zz_3               (_zz_3                           ), //i
    ._zz_4               (_zz_2_regNext                   )  //i
  );
  SingleKey singleKey_172 (
    .raw                 (_zz_73                          ), //i
    .filtered_valid      (singleKey_172_filtered_valid    ), //o
    .filtered_payload    (singleKey_172_filtered_payload  ), //o
    .CLK_50              (CLK_50                          ), //i
    ._zz_3               (_zz_3                           ), //i
    ._zz_4               (_zz_2_regNext                   )  //i
  );
  SingleKey singleKey_173 (
    .raw                 (_zz_74                          ), //i
    .filtered_valid      (singleKey_173_filtered_valid    ), //o
    .filtered_payload    (singleKey_173_filtered_payload  ), //o
    .CLK_50              (CLK_50                          ), //i
    ._zz_3               (_zz_3                           ), //i
    ._zz_4               (_zz_2_regNext                   )  //i
  );
  SingleKey singleKey_174 (
    .raw                 (_zz_75                          ), //i
    .filtered_valid      (singleKey_174_filtered_valid    ), //o
    .filtered_payload    (singleKey_174_filtered_payload  ), //o
    .CLK_50              (CLK_50                          ), //i
    ._zz_3               (_zz_3                           ), //i
    ._zz_4               (_zz_2_regNext                   )  //i
  );
  SingleKey singleKey_175 (
    .raw                 (_zz_76                          ), //i
    .filtered_valid      (singleKey_175_filtered_valid    ), //o
    .filtered_payload    (singleKey_175_filtered_payload  ), //o
    .CLK_50              (CLK_50                          ), //i
    ._zz_3               (_zz_3                           ), //i
    ._zz_4               (_zz_2_regNext                   )  //i
  );
  SingleKey singleKey_176 (
    .raw                 (_zz_77                          ), //i
    .filtered_valid      (singleKey_176_filtered_valid    ), //o
    .filtered_payload    (singleKey_176_filtered_payload  ), //o
    .CLK_50              (CLK_50                          ), //i
    ._zz_3               (_zz_3                           ), //i
    ._zz_4               (_zz_2_regNext                   )  //i
  );
  SingleKey singleKey_177 (
    .raw                 (_zz_78                          ), //i
    .filtered_valid      (singleKey_177_filtered_valid    ), //o
    .filtered_payload    (singleKey_177_filtered_payload  ), //o
    .CLK_50              (CLK_50                          ), //i
    ._zz_3               (_zz_3                           ), //i
    ._zz_4               (_zz_2_regNext                   )  //i
  );
  SingleKey singleKey_178 (
    .raw                 (_zz_79                          ), //i
    .filtered_valid      (singleKey_178_filtered_valid    ), //o
    .filtered_payload    (singleKey_178_filtered_payload  ), //o
    .CLK_50              (CLK_50                          ), //i
    ._zz_3               (_zz_3                           ), //i
    ._zz_4               (_zz_2_regNext                   )  //i
  );
  SingleKey singleKey_179 (
    .raw                 (_zz_80                          ), //i
    .filtered_valid      (singleKey_179_filtered_valid    ), //o
    .filtered_payload    (singleKey_179_filtered_payload  ), //o
    .CLK_50              (CLK_50                          ), //i
    ._zz_3               (_zz_3                           ), //i
    ._zz_4               (_zz_2_regNext                   )  //i
  );
  SingleKey singleKey_180 (
    .raw                 (_zz_81                          ), //i
    .filtered_valid      (singleKey_180_filtered_valid    ), //o
    .filtered_payload    (singleKey_180_filtered_payload  ), //o
    .CLK_50              (CLK_50                          ), //i
    ._zz_3               (_zz_3                           ), //i
    ._zz_4               (_zz_2_regNext                   )  //i
  );
  SingleKey singleKey_181 (
    .raw                 (_zz_82                          ), //i
    .filtered_valid      (singleKey_181_filtered_valid    ), //o
    .filtered_payload    (singleKey_181_filtered_payload  ), //o
    .CLK_50              (CLK_50                          ), //i
    ._zz_3               (_zz_3                           ), //i
    ._zz_4               (_zz_2_regNext                   )  //i
  );
  SingleKey singleKey_182 (
    .raw                 (_zz_83                          ), //i
    .filtered_valid      (singleKey_182_filtered_valid    ), //o
    .filtered_payload    (singleKey_182_filtered_payload  ), //o
    .CLK_50              (CLK_50                          ), //i
    ._zz_3               (_zz_3                           ), //i
    ._zz_4               (_zz_2_regNext                   )  //i
  );
  SingleKey singleKey_183 (
    .raw                 (_zz_84                          ), //i
    .filtered_valid      (singleKey_183_filtered_valid    ), //o
    .filtered_payload    (singleKey_183_filtered_payload  ), //o
    .CLK_50              (CLK_50                          ), //i
    ._zz_3               (_zz_3                           ), //i
    ._zz_4               (_zz_2_regNext                   )  //i
  );
  SingleKey singleKey_184 (
    .raw                 (_zz_85                          ), //i
    .filtered_valid      (singleKey_184_filtered_valid    ), //o
    .filtered_payload    (singleKey_184_filtered_payload  ), //o
    .CLK_50              (CLK_50                          ), //i
    ._zz_3               (_zz_3                           ), //i
    ._zz_4               (_zz_2_regNext                   )  //i
  );
  SingleKey singleKey_185 (
    .raw                 (_zz_86                          ), //i
    .filtered_valid      (singleKey_185_filtered_valid    ), //o
    .filtered_payload    (singleKey_185_filtered_payload  ), //o
    .CLK_50              (CLK_50                          ), //i
    ._zz_3               (_zz_3                           ), //i
    ._zz_4               (_zz_2_regNext                   )  //i
  );
  SingleKey singleKey_186 (
    .raw                 (_zz_87                          ), //i
    .filtered_valid      (singleKey_186_filtered_valid    ), //o
    .filtered_payload    (singleKey_186_filtered_payload  ), //o
    .CLK_50              (CLK_50                          ), //i
    ._zz_3               (_zz_3                           ), //i
    ._zz_4               (_zz_2_regNext                   )  //i
  );
  SingleKey singleKey_187 (
    .raw                 (_zz_88                          ), //i
    .filtered_valid      (singleKey_187_filtered_valid    ), //o
    .filtered_payload    (singleKey_187_filtered_payload  ), //o
    .CLK_50              (CLK_50                          ), //i
    ._zz_3               (_zz_3                           ), //i
    ._zz_4               (_zz_2_regNext                   )  //i
  );
  SingleKey singleKey_188 (
    .raw                 (_zz_89                          ), //i
    .filtered_valid      (singleKey_188_filtered_valid    ), //o
    .filtered_payload    (singleKey_188_filtered_payload  ), //o
    .CLK_50              (CLK_50                          ), //i
    ._zz_3               (_zz_3                           ), //i
    ._zz_4               (_zz_2_regNext                   )  //i
  );
  SingleKey singleKey_189 (
    .raw                 (_zz_90                          ), //i
    .filtered_valid      (singleKey_189_filtered_valid    ), //o
    .filtered_payload    (singleKey_189_filtered_payload  ), //o
    .CLK_50              (CLK_50                          ), //i
    ._zz_3               (_zz_3                           ), //i
    ._zz_4               (_zz_2_regNext                   )  //i
  );
  SingleKey singleKey_190 (
    .raw                 (_zz_91                          ), //i
    .filtered_valid      (singleKey_190_filtered_valid    ), //o
    .filtered_payload    (singleKey_190_filtered_payload  ), //o
    .CLK_50              (CLK_50                          ), //i
    ._zz_3               (_zz_3                           ), //i
    ._zz_4               (_zz_2_regNext                   )  //i
  );
  SingleKey singleKey_191 (
    .raw                 (_zz_92                          ), //i
    .filtered_valid      (singleKey_191_filtered_valid    ), //o
    .filtered_payload    (singleKey_191_filtered_payload  ), //o
    .CLK_50              (CLK_50                          ), //i
    ._zz_3               (_zz_3                           ), //i
    ._zz_4               (_zz_2_regNext                   )  //i
  );
  SingleKey singleKey_192 (
    .raw                 (_zz_93                          ), //i
    .filtered_valid      (singleKey_192_filtered_valid    ), //o
    .filtered_payload    (singleKey_192_filtered_payload  ), //o
    .CLK_50              (CLK_50                          ), //i
    ._zz_3               (_zz_3                           ), //i
    ._zz_4               (_zz_2_regNext                   )  //i
  );
  SingleKey singleKey_193 (
    .raw                 (_zz_94                          ), //i
    .filtered_valid      (singleKey_193_filtered_valid    ), //o
    .filtered_payload    (singleKey_193_filtered_payload  ), //o
    .CLK_50              (CLK_50                          ), //i
    ._zz_3               (_zz_3                           ), //i
    ._zz_4               (_zz_2_regNext                   )  //i
  );
  SingleKey singleKey_194 (
    .raw                 (_zz_95                          ), //i
    .filtered_valid      (singleKey_194_filtered_valid    ), //o
    .filtered_payload    (singleKey_194_filtered_payload  ), //o
    .CLK_50              (CLK_50                          ), //i
    ._zz_3               (_zz_3                           ), //i
    ._zz_4               (_zz_2_regNext                   )  //i
  );
  SingleKey singleKey_195 (
    .raw                 (_zz_96                          ), //i
    .filtered_valid      (singleKey_195_filtered_valid    ), //o
    .filtered_payload    (singleKey_195_filtered_payload  ), //o
    .CLK_50              (CLK_50                          ), //i
    ._zz_3               (_zz_3                           ), //i
    ._zz_4               (_zz_2_regNext                   )  //i
  );
  SingleKey singleKey_196 (
    .raw                 (_zz_97                          ), //i
    .filtered_valid      (singleKey_196_filtered_valid    ), //o
    .filtered_payload    (singleKey_196_filtered_payload  ), //o
    .CLK_50              (CLK_50                          ), //i
    ._zz_3               (_zz_3                           ), //i
    ._zz_4               (_zz_2_regNext                   )  //i
  );
  SingleKey singleKey_197 (
    .raw                 (_zz_98                          ), //i
    .filtered_valid      (singleKey_197_filtered_valid    ), //o
    .filtered_payload    (singleKey_197_filtered_payload  ), //o
    .CLK_50              (CLK_50                          ), //i
    ._zz_3               (_zz_3                           ), //i
    ._zz_4               (_zz_2_regNext                   )  //i
  );
  SingleKey singleKey_198 (
    .raw                 (_zz_99                          ), //i
    .filtered_valid      (singleKey_198_filtered_valid    ), //o
    .filtered_payload    (singleKey_198_filtered_payload  ), //o
    .CLK_50              (CLK_50                          ), //i
    ._zz_3               (_zz_3                           ), //i
    ._zz_4               (_zz_2_regNext                   )  //i
  );
  SingleKey singleKey_199 (
    .raw                 (_zz_100                         ), //i
    .filtered_valid      (singleKey_199_filtered_valid    ), //o
    .filtered_payload    (singleKey_199_filtered_payload  ), //o
    .CLK_50              (CLK_50                          ), //i
    ._zz_3               (_zz_3                           ), //i
    ._zz_4               (_zz_2_regNext                   )  //i
  );
  SingleKey singleKey_200 (
    .raw                 (_zz_101                         ), //i
    .filtered_valid      (singleKey_200_filtered_valid    ), //o
    .filtered_payload    (singleKey_200_filtered_payload  ), //o
    .CLK_50              (CLK_50                          ), //i
    ._zz_3               (_zz_3                           ), //i
    ._zz_4               (_zz_2_regNext                   )  //i
  );
  SingleKey singleKey_201 (
    .raw                 (_zz_102                         ), //i
    .filtered_valid      (singleKey_201_filtered_valid    ), //o
    .filtered_payload    (singleKey_201_filtered_payload  ), //o
    .CLK_50              (CLK_50                          ), //i
    ._zz_3               (_zz_3                           ), //i
    ._zz_4               (_zz_2_regNext                   )  //i
  );
  SingleKey singleKey_202 (
    .raw                 (_zz_103                         ), //i
    .filtered_valid      (singleKey_202_filtered_valid    ), //o
    .filtered_payload    (singleKey_202_filtered_payload  ), //o
    .CLK_50              (CLK_50                          ), //i
    ._zz_3               (_zz_3                           ), //i
    ._zz_4               (_zz_2_regNext                   )  //i
  );
  SingleKey singleKey_203 (
    .raw                 (_zz_104                         ), //i
    .filtered_valid      (singleKey_203_filtered_valid    ), //o
    .filtered_payload    (singleKey_203_filtered_payload  ), //o
    .CLK_50              (CLK_50                          ), //i
    ._zz_3               (_zz_3                           ), //i
    ._zz_4               (_zz_2_regNext                   )  //i
  );
  SingleKey singleKey_204 (
    .raw                 (_zz_105                         ), //i
    .filtered_valid      (singleKey_204_filtered_valid    ), //o
    .filtered_payload    (singleKey_204_filtered_payload  ), //o
    .CLK_50              (CLK_50                          ), //i
    ._zz_3               (_zz_3                           ), //i
    ._zz_4               (_zz_2_regNext                   )  //i
  );
  SingleKey singleKey_205 (
    .raw                 (_zz_106                         ), //i
    .filtered_valid      (singleKey_205_filtered_valid    ), //o
    .filtered_payload    (singleKey_205_filtered_payload  ), //o
    .CLK_50              (CLK_50                          ), //i
    ._zz_3               (_zz_3                           ), //i
    ._zz_4               (_zz_2_regNext                   )  //i
  );
  assign _zz_2 = (_zz_1 == 14'h270f);
  assign _zz_4 = key_down[0];
  assign keyStatus_0_valid = singleKey_103_filtered_valid;
  assign keyStatus_0_payload = singleKey_103_filtered_payload;
  assign _zz_5 = key_down[1];
  assign keyStatus_1_valid = singleKey_104_filtered_valid;
  assign keyStatus_1_payload = singleKey_104_filtered_payload;
  assign _zz_6 = key_down[2];
  assign keyStatus_2_valid = singleKey_105_filtered_valid;
  assign keyStatus_2_payload = singleKey_105_filtered_payload;
  assign _zz_7 = key_down[3];
  assign keyStatus_3_valid = singleKey_106_filtered_valid;
  assign keyStatus_3_payload = singleKey_106_filtered_payload;
  assign _zz_8 = key_down[4];
  assign keyStatus_4_valid = singleKey_107_filtered_valid;
  assign keyStatus_4_payload = singleKey_107_filtered_payload;
  assign _zz_9 = key_down[5];
  assign keyStatus_5_valid = singleKey_108_filtered_valid;
  assign keyStatus_5_payload = singleKey_108_filtered_payload;
  assign _zz_10 = key_down[6];
  assign keyStatus_6_valid = singleKey_109_filtered_valid;
  assign keyStatus_6_payload = singleKey_109_filtered_payload;
  assign _zz_11 = key_down[7];
  assign keyStatus_7_valid = singleKey_110_filtered_valid;
  assign keyStatus_7_payload = singleKey_110_filtered_payload;
  assign _zz_12 = key_down[8];
  assign keyStatus_8_valid = singleKey_111_filtered_valid;
  assign keyStatus_8_payload = singleKey_111_filtered_payload;
  assign _zz_13 = key_down[9];
  assign keyStatus_9_valid = singleKey_112_filtered_valid;
  assign keyStatus_9_payload = singleKey_112_filtered_payload;
  assign _zz_14 = key_down[10];
  assign keyStatus_10_valid = singleKey_113_filtered_valid;
  assign keyStatus_10_payload = singleKey_113_filtered_payload;
  assign _zz_15 = key_down[11];
  assign keyStatus_11_valid = singleKey_114_filtered_valid;
  assign keyStatus_11_payload = singleKey_114_filtered_payload;
  assign _zz_16 = key_down[12];
  assign keyStatus_12_valid = singleKey_115_filtered_valid;
  assign keyStatus_12_payload = singleKey_115_filtered_payload;
  assign _zz_17 = key_down[13];
  assign keyStatus_13_valid = singleKey_116_filtered_valid;
  assign keyStatus_13_payload = singleKey_116_filtered_payload;
  assign _zz_18 = key_down[14];
  assign keyStatus_14_valid = singleKey_117_filtered_valid;
  assign keyStatus_14_payload = singleKey_117_filtered_payload;
  assign _zz_19 = key_down[15];
  assign keyStatus_15_valid = singleKey_118_filtered_valid;
  assign keyStatus_15_payload = singleKey_118_filtered_payload;
  assign _zz_20 = key_down[16];
  assign keyStatus_16_valid = singleKey_119_filtered_valid;
  assign keyStatus_16_payload = singleKey_119_filtered_payload;
  assign _zz_21 = key_down[17];
  assign keyStatus_17_valid = singleKey_120_filtered_valid;
  assign keyStatus_17_payload = singleKey_120_filtered_payload;
  assign _zz_22 = key_down[18];
  assign keyStatus_18_valid = singleKey_121_filtered_valid;
  assign keyStatus_18_payload = singleKey_121_filtered_payload;
  assign _zz_23 = key_down[19];
  assign keyStatus_19_valid = singleKey_122_filtered_valid;
  assign keyStatus_19_payload = singleKey_122_filtered_payload;
  assign _zz_24 = key_down[20];
  assign keyStatus_20_valid = singleKey_123_filtered_valid;
  assign keyStatus_20_payload = singleKey_123_filtered_payload;
  assign _zz_25 = key_down[21];
  assign keyStatus_21_valid = singleKey_124_filtered_valid;
  assign keyStatus_21_payload = singleKey_124_filtered_payload;
  assign _zz_26 = key_down[22];
  assign keyStatus_22_valid = singleKey_125_filtered_valid;
  assign keyStatus_22_payload = singleKey_125_filtered_payload;
  assign _zz_27 = key_down[23];
  assign keyStatus_23_valid = singleKey_126_filtered_valid;
  assign keyStatus_23_payload = singleKey_126_filtered_payload;
  assign _zz_28 = key_down[24];
  assign keyStatus_24_valid = singleKey_127_filtered_valid;
  assign keyStatus_24_payload = singleKey_127_filtered_payload;
  assign _zz_29 = key_down[25];
  assign keyStatus_25_valid = singleKey_128_filtered_valid;
  assign keyStatus_25_payload = singleKey_128_filtered_payload;
  assign _zz_30 = key_down[26];
  assign keyStatus_26_valid = singleKey_129_filtered_valid;
  assign keyStatus_26_payload = singleKey_129_filtered_payload;
  assign _zz_31 = key_down[27];
  assign keyStatus_27_valid = singleKey_130_filtered_valid;
  assign keyStatus_27_payload = singleKey_130_filtered_payload;
  assign _zz_32 = key_down[28];
  assign keyStatus_28_valid = singleKey_131_filtered_valid;
  assign keyStatus_28_payload = singleKey_131_filtered_payload;
  assign _zz_33 = key_down[29];
  assign keyStatus_29_valid = singleKey_132_filtered_valid;
  assign keyStatus_29_payload = singleKey_132_filtered_payload;
  assign _zz_34 = key_down[30];
  assign keyStatus_30_valid = singleKey_133_filtered_valid;
  assign keyStatus_30_payload = singleKey_133_filtered_payload;
  assign _zz_35 = key_down[31];
  assign keyStatus_31_valid = singleKey_134_filtered_valid;
  assign keyStatus_31_payload = singleKey_134_filtered_payload;
  assign _zz_36 = key_down[32];
  assign keyStatus_32_valid = singleKey_135_filtered_valid;
  assign keyStatus_32_payload = singleKey_135_filtered_payload;
  assign _zz_37 = key_down[33];
  assign keyStatus_33_valid = singleKey_136_filtered_valid;
  assign keyStatus_33_payload = singleKey_136_filtered_payload;
  assign _zz_38 = key_down[34];
  assign keyStatus_34_valid = singleKey_137_filtered_valid;
  assign keyStatus_34_payload = singleKey_137_filtered_payload;
  assign _zz_39 = key_down[35];
  assign keyStatus_35_valid = singleKey_138_filtered_valid;
  assign keyStatus_35_payload = singleKey_138_filtered_payload;
  assign _zz_40 = key_down[36];
  assign keyStatus_36_valid = singleKey_139_filtered_valid;
  assign keyStatus_36_payload = singleKey_139_filtered_payload;
  assign _zz_41 = key_down[37];
  assign keyStatus_37_valid = singleKey_140_filtered_valid;
  assign keyStatus_37_payload = singleKey_140_filtered_payload;
  assign _zz_42 = key_down[38];
  assign keyStatus_38_valid = singleKey_141_filtered_valid;
  assign keyStatus_38_payload = singleKey_141_filtered_payload;
  assign _zz_43 = key_down[39];
  assign keyStatus_39_valid = singleKey_142_filtered_valid;
  assign keyStatus_39_payload = singleKey_142_filtered_payload;
  assign _zz_44 = key_down[40];
  assign keyStatus_40_valid = singleKey_143_filtered_valid;
  assign keyStatus_40_payload = singleKey_143_filtered_payload;
  assign _zz_45 = key_down[41];
  assign keyStatus_41_valid = singleKey_144_filtered_valid;
  assign keyStatus_41_payload = singleKey_144_filtered_payload;
  assign _zz_46 = key_down[42];
  assign keyStatus_42_valid = singleKey_145_filtered_valid;
  assign keyStatus_42_payload = singleKey_145_filtered_payload;
  assign _zz_47 = key_down[43];
  assign keyStatus_43_valid = singleKey_146_filtered_valid;
  assign keyStatus_43_payload = singleKey_146_filtered_payload;
  assign _zz_48 = key_down[44];
  assign keyStatus_44_valid = singleKey_147_filtered_valid;
  assign keyStatus_44_payload = singleKey_147_filtered_payload;
  assign _zz_49 = key_down[45];
  assign keyStatus_45_valid = singleKey_148_filtered_valid;
  assign keyStatus_45_payload = singleKey_148_filtered_payload;
  assign _zz_50 = key_down[46];
  assign keyStatus_46_valid = singleKey_149_filtered_valid;
  assign keyStatus_46_payload = singleKey_149_filtered_payload;
  assign _zz_51 = key_down[47];
  assign keyStatus_47_valid = singleKey_150_filtered_valid;
  assign keyStatus_47_payload = singleKey_150_filtered_payload;
  assign _zz_52 = key_down[48];
  assign keyStatus_48_valid = singleKey_151_filtered_valid;
  assign keyStatus_48_payload = singleKey_151_filtered_payload;
  assign _zz_53 = key_down[49];
  assign keyStatus_49_valid = singleKey_152_filtered_valid;
  assign keyStatus_49_payload = singleKey_152_filtered_payload;
  assign _zz_54 = key_down[50];
  assign keyStatus_50_valid = singleKey_153_filtered_valid;
  assign keyStatus_50_payload = singleKey_153_filtered_payload;
  assign _zz_55 = key_down[51];
  assign keyStatus_51_valid = singleKey_154_filtered_valid;
  assign keyStatus_51_payload = singleKey_154_filtered_payload;
  assign _zz_56 = key_down[52];
  assign keyStatus_52_valid = singleKey_155_filtered_valid;
  assign keyStatus_52_payload = singleKey_155_filtered_payload;
  assign _zz_57 = key_down[53];
  assign keyStatus_53_valid = singleKey_156_filtered_valid;
  assign keyStatus_53_payload = singleKey_156_filtered_payload;
  assign _zz_58 = key_down[54];
  assign keyStatus_54_valid = singleKey_157_filtered_valid;
  assign keyStatus_54_payload = singleKey_157_filtered_payload;
  assign _zz_59 = key_down[55];
  assign keyStatus_55_valid = singleKey_158_filtered_valid;
  assign keyStatus_55_payload = singleKey_158_filtered_payload;
  assign _zz_60 = key_down[56];
  assign keyStatus_56_valid = singleKey_159_filtered_valid;
  assign keyStatus_56_payload = singleKey_159_filtered_payload;
  assign _zz_61 = key_down[57];
  assign keyStatus_57_valid = singleKey_160_filtered_valid;
  assign keyStatus_57_payload = singleKey_160_filtered_payload;
  assign _zz_62 = key_down[58];
  assign keyStatus_58_valid = singleKey_161_filtered_valid;
  assign keyStatus_58_payload = singleKey_161_filtered_payload;
  assign _zz_63 = key_down[59];
  assign keyStatus_59_valid = singleKey_162_filtered_valid;
  assign keyStatus_59_payload = singleKey_162_filtered_payload;
  assign _zz_64 = key_down[60];
  assign keyStatus_60_valid = singleKey_163_filtered_valid;
  assign keyStatus_60_payload = singleKey_163_filtered_payload;
  assign _zz_65 = key_down[61];
  assign keyStatus_61_valid = singleKey_164_filtered_valid;
  assign keyStatus_61_payload = singleKey_164_filtered_payload;
  assign _zz_66 = key_down[62];
  assign keyStatus_62_valid = singleKey_165_filtered_valid;
  assign keyStatus_62_payload = singleKey_165_filtered_payload;
  assign _zz_67 = key_down[63];
  assign keyStatus_63_valid = singleKey_166_filtered_valid;
  assign keyStatus_63_payload = singleKey_166_filtered_payload;
  assign _zz_68 = key_down[64];
  assign keyStatus_64_valid = singleKey_167_filtered_valid;
  assign keyStatus_64_payload = singleKey_167_filtered_payload;
  assign _zz_69 = key_down[65];
  assign keyStatus_65_valid = singleKey_168_filtered_valid;
  assign keyStatus_65_payload = singleKey_168_filtered_payload;
  assign _zz_70 = key_down[66];
  assign keyStatus_66_valid = singleKey_169_filtered_valid;
  assign keyStatus_66_payload = singleKey_169_filtered_payload;
  assign _zz_71 = key_down[67];
  assign keyStatus_67_valid = singleKey_170_filtered_valid;
  assign keyStatus_67_payload = singleKey_170_filtered_payload;
  assign _zz_72 = key_down[68];
  assign keyStatus_68_valid = singleKey_171_filtered_valid;
  assign keyStatus_68_payload = singleKey_171_filtered_payload;
  assign _zz_73 = key_down[69];
  assign keyStatus_69_valid = singleKey_172_filtered_valid;
  assign keyStatus_69_payload = singleKey_172_filtered_payload;
  assign _zz_74 = key_down[70];
  assign keyStatus_70_valid = singleKey_173_filtered_valid;
  assign keyStatus_70_payload = singleKey_173_filtered_payload;
  assign _zz_75 = key_down[71];
  assign keyStatus_71_valid = singleKey_174_filtered_valid;
  assign keyStatus_71_payload = singleKey_174_filtered_payload;
  assign _zz_76 = key_down[72];
  assign keyStatus_72_valid = singleKey_175_filtered_valid;
  assign keyStatus_72_payload = singleKey_175_filtered_payload;
  assign _zz_77 = key_down[73];
  assign keyStatus_73_valid = singleKey_176_filtered_valid;
  assign keyStatus_73_payload = singleKey_176_filtered_payload;
  assign _zz_78 = key_down[74];
  assign keyStatus_74_valid = singleKey_177_filtered_valid;
  assign keyStatus_74_payload = singleKey_177_filtered_payload;
  assign _zz_79 = key_down[75];
  assign keyStatus_75_valid = singleKey_178_filtered_valid;
  assign keyStatus_75_payload = singleKey_178_filtered_payload;
  assign _zz_80 = key_down[76];
  assign keyStatus_76_valid = singleKey_179_filtered_valid;
  assign keyStatus_76_payload = singleKey_179_filtered_payload;
  assign _zz_81 = key_down[77];
  assign keyStatus_77_valid = singleKey_180_filtered_valid;
  assign keyStatus_77_payload = singleKey_180_filtered_payload;
  assign _zz_82 = key_down[78];
  assign keyStatus_78_valid = singleKey_181_filtered_valid;
  assign keyStatus_78_payload = singleKey_181_filtered_payload;
  assign _zz_83 = key_down[79];
  assign keyStatus_79_valid = singleKey_182_filtered_valid;
  assign keyStatus_79_payload = singleKey_182_filtered_payload;
  assign _zz_84 = key_down[80];
  assign keyStatus_80_valid = singleKey_183_filtered_valid;
  assign keyStatus_80_payload = singleKey_183_filtered_payload;
  assign _zz_85 = key_down[81];
  assign keyStatus_81_valid = singleKey_184_filtered_valid;
  assign keyStatus_81_payload = singleKey_184_filtered_payload;
  assign _zz_86 = key_down[82];
  assign keyStatus_82_valid = singleKey_185_filtered_valid;
  assign keyStatus_82_payload = singleKey_185_filtered_payload;
  assign _zz_87 = key_down[83];
  assign keyStatus_83_valid = singleKey_186_filtered_valid;
  assign keyStatus_83_payload = singleKey_186_filtered_payload;
  assign _zz_88 = key_down[84];
  assign keyStatus_84_valid = singleKey_187_filtered_valid;
  assign keyStatus_84_payload = singleKey_187_filtered_payload;
  assign _zz_89 = key_down[85];
  assign keyStatus_85_valid = singleKey_188_filtered_valid;
  assign keyStatus_85_payload = singleKey_188_filtered_payload;
  assign _zz_90 = key_down[86];
  assign keyStatus_86_valid = singleKey_189_filtered_valid;
  assign keyStatus_86_payload = singleKey_189_filtered_payload;
  assign _zz_91 = key_down[87];
  assign keyStatus_87_valid = singleKey_190_filtered_valid;
  assign keyStatus_87_payload = singleKey_190_filtered_payload;
  assign _zz_92 = key_down[88];
  assign keyStatus_88_valid = singleKey_191_filtered_valid;
  assign keyStatus_88_payload = singleKey_191_filtered_payload;
  assign _zz_93 = key_down[89];
  assign keyStatus_89_valid = singleKey_192_filtered_valid;
  assign keyStatus_89_payload = singleKey_192_filtered_payload;
  assign _zz_94 = key_down[90];
  assign keyStatus_90_valid = singleKey_193_filtered_valid;
  assign keyStatus_90_payload = singleKey_193_filtered_payload;
  assign _zz_95 = key_down[91];
  assign keyStatus_91_valid = singleKey_194_filtered_valid;
  assign keyStatus_91_payload = singleKey_194_filtered_payload;
  assign _zz_96 = key_down[92];
  assign keyStatus_92_valid = singleKey_195_filtered_valid;
  assign keyStatus_92_payload = singleKey_195_filtered_payload;
  assign _zz_97 = key_down[93];
  assign keyStatus_93_valid = singleKey_196_filtered_valid;
  assign keyStatus_93_payload = singleKey_196_filtered_payload;
  assign _zz_98 = key_down[94];
  assign keyStatus_94_valid = singleKey_197_filtered_valid;
  assign keyStatus_94_payload = singleKey_197_filtered_payload;
  assign _zz_99 = key_down[95];
  assign keyStatus_95_valid = singleKey_198_filtered_valid;
  assign keyStatus_95_payload = singleKey_198_filtered_payload;
  assign _zz_100 = key_down[96];
  assign keyStatus_96_valid = singleKey_199_filtered_valid;
  assign keyStatus_96_payload = singleKey_199_filtered_payload;
  assign _zz_101 = key_down[97];
  assign keyStatus_97_valid = singleKey_200_filtered_valid;
  assign keyStatus_97_payload = singleKey_200_filtered_payload;
  assign _zz_102 = key_down[98];
  assign keyStatus_98_valid = singleKey_201_filtered_valid;
  assign keyStatus_98_payload = singleKey_201_filtered_payload;
  assign _zz_103 = key_down[99];
  assign keyStatus_99_valid = singleKey_202_filtered_valid;
  assign keyStatus_99_payload = singleKey_202_filtered_payload;
  assign _zz_104 = key_down[100];
  assign keyStatus_100_valid = singleKey_203_filtered_valid;
  assign keyStatus_100_payload = singleKey_203_filtered_payload;
  assign _zz_105 = key_down[101];
  assign keyStatus_101_valid = singleKey_204_filtered_valid;
  assign keyStatus_101_payload = singleKey_204_filtered_payload;
  assign _zz_106 = key_down[102];
  assign keyStatus_102_valid = singleKey_205_filtered_valid;
  assign keyStatus_102_payload = singleKey_205_filtered_payload;
  always @ (posedge CLK_50 or posedge _zz_3) begin
    if (_zz_3) begin
      _zz_1 <= 14'h0;
      _zz_2_regNext <= 1'b0;
    end else begin
      _zz_1 <= (_zz_1 + 14'h0001);
      if(_zz_2)begin
        _zz_1 <= 14'h0;
      end
      _zz_2_regNext <= _zz_2;
    end
  end


endmodule

module UartCtrlRx (
  input      [2:0]    io_configFrame_dataLength,
  input      `UartStopType_defaultEncoding_type io_configFrame_stop,
  input      `UartParityType_defaultEncoding_type io_configFrame_parity,
  input               io_samplingTick,
  output              io_read_valid,
  input               io_read_ready,
  output     [7:0]    io_read_payload,
  input               io_rxd,
  output              io_rts,
  output reg          io_error,
  output              io_break,
  input               CLK_50,
  input               _zz_2
);
  wire                io_rxd_buffercc_io_dataOut;
  wire                _zz_3;
  wire                _zz_4;
  wire                _zz_5;
  wire                _zz_6;
  wire       [0:0]    _zz_7;
  wire       [2:0]    _zz_8;
  wire                _zz_9;
  wire                _zz_10;
  wire                _zz_11;
  wire                _zz_12;
  wire                _zz_13;
  wire                _zz_14;
  wire                _zz_15;
  reg                 _zz_1;
  wire                sampler_synchroniser;
  wire                sampler_samples_0;
  reg                 sampler_samples_1;
  reg                 sampler_samples_2;
  reg                 sampler_samples_3;
  reg                 sampler_samples_4;
  reg                 sampler_value;
  reg                 sampler_tick;
  reg        [2:0]    bitTimer_counter;
  reg                 bitTimer_tick;
  reg        [2:0]    bitCounter_value;
  reg        [6:0]    break_counter;
  wire                break_valid;
  reg        `UartCtrlRxState_defaultEncoding_type stateMachine_state;
  reg                 stateMachine_parity;
  reg        [7:0]    stateMachine_shifter;
  reg                 stateMachine_validReg;
  `ifndef SYNTHESIS
  reg [23:0] io_configFrame_stop_string;
  reg [31:0] io_configFrame_parity_string;
  reg [47:0] stateMachine_state_string;
  `endif


  assign _zz_3 = (stateMachine_parity == sampler_value);
  assign _zz_4 = (! sampler_value);
  assign _zz_5 = ((sampler_tick && (! sampler_value)) && (! break_valid));
  assign _zz_6 = (bitCounter_value == io_configFrame_dataLength);
  assign _zz_7 = ((io_configFrame_stop == `UartStopType_defaultEncoding_ONE) ? 1'b0 : 1'b1);
  assign _zz_8 = {2'd0, _zz_7};
  assign _zz_9 = ((((1'b0 || ((_zz_14 && sampler_samples_1) && sampler_samples_2)) || (((_zz_15 && sampler_samples_0) && sampler_samples_1) && sampler_samples_3)) || (((1'b1 && sampler_samples_0) && sampler_samples_2) && sampler_samples_3)) || (((1'b1 && sampler_samples_1) && sampler_samples_2) && sampler_samples_3));
  assign _zz_10 = (((1'b1 && sampler_samples_0) && sampler_samples_1) && sampler_samples_4);
  assign _zz_11 = ((1'b1 && sampler_samples_0) && sampler_samples_2);
  assign _zz_12 = (1'b1 && sampler_samples_1);
  assign _zz_13 = 1'b1;
  assign _zz_14 = (1'b1 && sampler_samples_0);
  assign _zz_15 = 1'b1;
  BufferCC io_rxd_buffercc (
    .io_dataIn     (io_rxd                      ), //i
    .io_dataOut    (io_rxd_buffercc_io_dataOut  ), //o
    .CLK_50        (CLK_50                      ), //i
    ._zz_1         (_zz_2                       )  //i
  );
  `ifndef SYNTHESIS
  always @(*) begin
    case(io_configFrame_stop)
      `UartStopType_defaultEncoding_ONE : io_configFrame_stop_string = "ONE";
      `UartStopType_defaultEncoding_TWO : io_configFrame_stop_string = "TWO";
      default : io_configFrame_stop_string = "???";
    endcase
  end
  always @(*) begin
    case(io_configFrame_parity)
      `UartParityType_defaultEncoding_NONE : io_configFrame_parity_string = "NONE";
      `UartParityType_defaultEncoding_EVEN : io_configFrame_parity_string = "EVEN";
      `UartParityType_defaultEncoding_ODD : io_configFrame_parity_string = "ODD ";
      default : io_configFrame_parity_string = "????";
    endcase
  end
  always @(*) begin
    case(stateMachine_state)
      `UartCtrlRxState_defaultEncoding_IDLE : stateMachine_state_string = "IDLE  ";
      `UartCtrlRxState_defaultEncoding_START : stateMachine_state_string = "START ";
      `UartCtrlRxState_defaultEncoding_DATA : stateMachine_state_string = "DATA  ";
      `UartCtrlRxState_defaultEncoding_PARITY : stateMachine_state_string = "PARITY";
      `UartCtrlRxState_defaultEncoding_STOP : stateMachine_state_string = "STOP  ";
      default : stateMachine_state_string = "??????";
    endcase
  end
  `endif

  always @ (*) begin
    io_error = 1'b0;
    case(stateMachine_state)
      `UartCtrlRxState_defaultEncoding_IDLE : begin
      end
      `UartCtrlRxState_defaultEncoding_START : begin
      end
      `UartCtrlRxState_defaultEncoding_DATA : begin
      end
      `UartCtrlRxState_defaultEncoding_PARITY : begin
        if(bitTimer_tick)begin
          if(! _zz_3) begin
            io_error = 1'b1;
          end
        end
      end
      default : begin
        if(bitTimer_tick)begin
          if(_zz_4)begin
            io_error = 1'b1;
          end
        end
      end
    endcase
  end

  assign io_rts = _zz_1;
  assign sampler_synchroniser = io_rxd_buffercc_io_dataOut;
  assign sampler_samples_0 = sampler_synchroniser;
  always @ (*) begin
    bitTimer_tick = 1'b0;
    if(sampler_tick)begin
      if((bitTimer_counter == 3'b000))begin
        bitTimer_tick = 1'b1;
      end
    end
  end

  assign break_valid = (break_counter == 7'h68);
  assign io_break = break_valid;
  assign io_read_valid = stateMachine_validReg;
  assign io_read_payload = stateMachine_shifter;
  always @ (posedge CLK_50 or posedge _zz_2) begin
    if (_zz_2) begin
      _zz_1 <= 1'b0;
      sampler_samples_1 <= 1'b1;
      sampler_samples_2 <= 1'b1;
      sampler_samples_3 <= 1'b1;
      sampler_samples_4 <= 1'b1;
      sampler_value <= 1'b1;
      sampler_tick <= 1'b0;
      break_counter <= 7'h0;
      stateMachine_state <= `UartCtrlRxState_defaultEncoding_IDLE;
      stateMachine_validReg <= 1'b0;
    end else begin
      _zz_1 <= (! io_read_ready);
      if(io_samplingTick)begin
        sampler_samples_1 <= sampler_samples_0;
      end
      if(io_samplingTick)begin
        sampler_samples_2 <= sampler_samples_1;
      end
      if(io_samplingTick)begin
        sampler_samples_3 <= sampler_samples_2;
      end
      if(io_samplingTick)begin
        sampler_samples_4 <= sampler_samples_3;
      end
      sampler_value <= ((((((_zz_9 || _zz_10) || (_zz_11 && sampler_samples_4)) || ((_zz_12 && sampler_samples_2) && sampler_samples_4)) || (((_zz_13 && sampler_samples_0) && sampler_samples_3) && sampler_samples_4)) || (((1'b1 && sampler_samples_1) && sampler_samples_3) && sampler_samples_4)) || (((1'b1 && sampler_samples_2) && sampler_samples_3) && sampler_samples_4));
      sampler_tick <= io_samplingTick;
      if(sampler_value)begin
        break_counter <= 7'h0;
      end else begin
        if((io_samplingTick && (! break_valid)))begin
          break_counter <= (break_counter + 7'h01);
        end
      end
      stateMachine_validReg <= 1'b0;
      case(stateMachine_state)
        `UartCtrlRxState_defaultEncoding_IDLE : begin
          if(_zz_5)begin
            stateMachine_state <= `UartCtrlRxState_defaultEncoding_START;
          end
        end
        `UartCtrlRxState_defaultEncoding_START : begin
          if(bitTimer_tick)begin
            stateMachine_state <= `UartCtrlRxState_defaultEncoding_DATA;
            if((sampler_value == 1'b1))begin
              stateMachine_state <= `UartCtrlRxState_defaultEncoding_IDLE;
            end
          end
        end
        `UartCtrlRxState_defaultEncoding_DATA : begin
          if(bitTimer_tick)begin
            if(_zz_6)begin
              if((io_configFrame_parity == `UartParityType_defaultEncoding_NONE))begin
                stateMachine_state <= `UartCtrlRxState_defaultEncoding_STOP;
                stateMachine_validReg <= 1'b1;
              end else begin
                stateMachine_state <= `UartCtrlRxState_defaultEncoding_PARITY;
              end
            end
          end
        end
        `UartCtrlRxState_defaultEncoding_PARITY : begin
          if(bitTimer_tick)begin
            if(_zz_3)begin
              stateMachine_state <= `UartCtrlRxState_defaultEncoding_STOP;
              stateMachine_validReg <= 1'b1;
            end else begin
              stateMachine_state <= `UartCtrlRxState_defaultEncoding_IDLE;
            end
          end
        end
        default : begin
          if(bitTimer_tick)begin
            if(_zz_4)begin
              stateMachine_state <= `UartCtrlRxState_defaultEncoding_IDLE;
            end else begin
              if((bitCounter_value == _zz_8))begin
                stateMachine_state <= `UartCtrlRxState_defaultEncoding_IDLE;
              end
            end
          end
        end
      endcase
    end
  end

  always @ (posedge CLK_50) begin
    if(sampler_tick)begin
      bitTimer_counter <= (bitTimer_counter - 3'b001);
    end
    if(bitTimer_tick)begin
      bitCounter_value <= (bitCounter_value + 3'b001);
    end
    if(bitTimer_tick)begin
      stateMachine_parity <= (stateMachine_parity ^ sampler_value);
    end
    case(stateMachine_state)
      `UartCtrlRxState_defaultEncoding_IDLE : begin
        if(_zz_5)begin
          bitTimer_counter <= 3'b010;
        end
      end
      `UartCtrlRxState_defaultEncoding_START : begin
        if(bitTimer_tick)begin
          bitCounter_value <= 3'b000;
          stateMachine_parity <= (io_configFrame_parity == `UartParityType_defaultEncoding_ODD);
        end
      end
      `UartCtrlRxState_defaultEncoding_DATA : begin
        if(bitTimer_tick)begin
          stateMachine_shifter[bitCounter_value] <= sampler_value;
          if(_zz_6)begin
            bitCounter_value <= 3'b000;
          end
        end
      end
      `UartCtrlRxState_defaultEncoding_PARITY : begin
        if(bitTimer_tick)begin
          bitCounter_value <= 3'b000;
        end
      end
      default : begin
      end
    endcase
  end


endmodule

module UartCtrlTx (
  input      [2:0]    io_configFrame_dataLength,
  input      `UartStopType_defaultEncoding_type io_configFrame_stop,
  input      `UartParityType_defaultEncoding_type io_configFrame_parity,
  input               io_samplingTick,
  input               io_write_valid,
  output reg          io_write_ready,
  input      [7:0]    io_write_payload,
  input               io_cts,
  output              io_txd,
  input               io_break,
  input               CLK_50,
  input               _zz_2
);
  wire                _zz_3;
  wire       [0:0]    _zz_4;
  wire       [2:0]    _zz_5;
  wire       [0:0]    _zz_6;
  wire       [2:0]    _zz_7;
  reg                 clockDivider_counter_willIncrement;
  wire                clockDivider_counter_willClear;
  reg        [2:0]    clockDivider_counter_valueNext;
  reg        [2:0]    clockDivider_counter_value;
  wire                clockDivider_counter_willOverflowIfInc;
  wire                clockDivider_counter_willOverflow;
  reg        [2:0]    tickCounter_value;
  reg        `UartCtrlTxState_defaultEncoding_type stateMachine_state;
  reg                 stateMachine_parity;
  reg                 stateMachine_txd;
  reg                 _zz_1;
  `ifndef SYNTHESIS
  reg [23:0] io_configFrame_stop_string;
  reg [31:0] io_configFrame_parity_string;
  reg [47:0] stateMachine_state_string;
  `endif


  assign _zz_3 = (tickCounter_value == io_configFrame_dataLength);
  assign _zz_4 = clockDivider_counter_willIncrement;
  assign _zz_5 = {2'd0, _zz_4};
  assign _zz_6 = ((io_configFrame_stop == `UartStopType_defaultEncoding_ONE) ? 1'b0 : 1'b1);
  assign _zz_7 = {2'd0, _zz_6};
  `ifndef SYNTHESIS
  always @(*) begin
    case(io_configFrame_stop)
      `UartStopType_defaultEncoding_ONE : io_configFrame_stop_string = "ONE";
      `UartStopType_defaultEncoding_TWO : io_configFrame_stop_string = "TWO";
      default : io_configFrame_stop_string = "???";
    endcase
  end
  always @(*) begin
    case(io_configFrame_parity)
      `UartParityType_defaultEncoding_NONE : io_configFrame_parity_string = "NONE";
      `UartParityType_defaultEncoding_EVEN : io_configFrame_parity_string = "EVEN";
      `UartParityType_defaultEncoding_ODD : io_configFrame_parity_string = "ODD ";
      default : io_configFrame_parity_string = "????";
    endcase
  end
  always @(*) begin
    case(stateMachine_state)
      `UartCtrlTxState_defaultEncoding_IDLE : stateMachine_state_string = "IDLE  ";
      `UartCtrlTxState_defaultEncoding_START : stateMachine_state_string = "START ";
      `UartCtrlTxState_defaultEncoding_DATA : stateMachine_state_string = "DATA  ";
      `UartCtrlTxState_defaultEncoding_PARITY : stateMachine_state_string = "PARITY";
      `UartCtrlTxState_defaultEncoding_STOP : stateMachine_state_string = "STOP  ";
      default : stateMachine_state_string = "??????";
    endcase
  end
  `endif

  always @ (*) begin
    clockDivider_counter_willIncrement = 1'b0;
    if(io_samplingTick)begin
      clockDivider_counter_willIncrement = 1'b1;
    end
  end

  assign clockDivider_counter_willClear = 1'b0;
  assign clockDivider_counter_willOverflowIfInc = (clockDivider_counter_value == 3'b111);
  assign clockDivider_counter_willOverflow = (clockDivider_counter_willOverflowIfInc && clockDivider_counter_willIncrement);
  always @ (*) begin
    clockDivider_counter_valueNext = (clockDivider_counter_value + _zz_5);
    if(clockDivider_counter_willClear)begin
      clockDivider_counter_valueNext = 3'b000;
    end
  end

  always @ (*) begin
    stateMachine_txd = 1'b1;
    case(stateMachine_state)
      `UartCtrlTxState_defaultEncoding_IDLE : begin
      end
      `UartCtrlTxState_defaultEncoding_START : begin
        stateMachine_txd = 1'b0;
      end
      `UartCtrlTxState_defaultEncoding_DATA : begin
        stateMachine_txd = io_write_payload[tickCounter_value];
      end
      `UartCtrlTxState_defaultEncoding_PARITY : begin
        stateMachine_txd = stateMachine_parity;
      end
      default : begin
      end
    endcase
  end

  always @ (*) begin
    io_write_ready = io_break;
    case(stateMachine_state)
      `UartCtrlTxState_defaultEncoding_IDLE : begin
      end
      `UartCtrlTxState_defaultEncoding_START : begin
      end
      `UartCtrlTxState_defaultEncoding_DATA : begin
        if(clockDivider_counter_willOverflow)begin
          if(_zz_3)begin
            io_write_ready = 1'b1;
          end
        end
      end
      `UartCtrlTxState_defaultEncoding_PARITY : begin
      end
      default : begin
      end
    endcase
  end

  assign io_txd = _zz_1;
  always @ (posedge CLK_50 or posedge _zz_2) begin
    if (_zz_2) begin
      clockDivider_counter_value <= 3'b000;
      stateMachine_state <= `UartCtrlTxState_defaultEncoding_IDLE;
      _zz_1 <= 1'b1;
    end else begin
      clockDivider_counter_value <= clockDivider_counter_valueNext;
      case(stateMachine_state)
        `UartCtrlTxState_defaultEncoding_IDLE : begin
          if(((io_write_valid && (! io_cts)) && clockDivider_counter_willOverflow))begin
            stateMachine_state <= `UartCtrlTxState_defaultEncoding_START;
          end
        end
        `UartCtrlTxState_defaultEncoding_START : begin
          if(clockDivider_counter_willOverflow)begin
            stateMachine_state <= `UartCtrlTxState_defaultEncoding_DATA;
          end
        end
        `UartCtrlTxState_defaultEncoding_DATA : begin
          if(clockDivider_counter_willOverflow)begin
            if(_zz_3)begin
              if((io_configFrame_parity == `UartParityType_defaultEncoding_NONE))begin
                stateMachine_state <= `UartCtrlTxState_defaultEncoding_STOP;
              end else begin
                stateMachine_state <= `UartCtrlTxState_defaultEncoding_PARITY;
              end
            end
          end
        end
        `UartCtrlTxState_defaultEncoding_PARITY : begin
          if(clockDivider_counter_willOverflow)begin
            stateMachine_state <= `UartCtrlTxState_defaultEncoding_STOP;
          end
        end
        default : begin
          if(clockDivider_counter_willOverflow)begin
            if((tickCounter_value == _zz_7))begin
              stateMachine_state <= (io_write_valid ? `UartCtrlTxState_defaultEncoding_START : `UartCtrlTxState_defaultEncoding_IDLE);
            end
          end
        end
      endcase
      _zz_1 <= (stateMachine_txd && (! io_break));
    end
  end

  always @ (posedge CLK_50) begin
    if(clockDivider_counter_willOverflow)begin
      tickCounter_value <= (tickCounter_value + 3'b001);
    end
    if(clockDivider_counter_willOverflow)begin
      stateMachine_parity <= (stateMachine_parity ^ stateMachine_txd);
    end
    case(stateMachine_state)
      `UartCtrlTxState_defaultEncoding_IDLE : begin
      end
      `UartCtrlTxState_defaultEncoding_START : begin
        if(clockDivider_counter_willOverflow)begin
          stateMachine_parity <= (io_configFrame_parity == `UartParityType_defaultEncoding_ODD);
          tickCounter_value <= 3'b000;
        end
      end
      `UartCtrlTxState_defaultEncoding_DATA : begin
        if(clockDivider_counter_willOverflow)begin
          if(_zz_3)begin
            tickCounter_value <= 3'b000;
          end
        end
      end
      `UartCtrlTxState_defaultEncoding_PARITY : begin
        if(clockDivider_counter_willOverflow)begin
          tickCounter_value <= 3'b000;
        end
      end
      default : begin
      end
    endcase
  end


endmodule

//SingleKey replaced by SingleKey

//SingleKey replaced by SingleKey

//SingleKey replaced by SingleKey

//SingleKey replaced by SingleKey

//SingleKey replaced by SingleKey

//SingleKey replaced by SingleKey

//SingleKey replaced by SingleKey

//SingleKey replaced by SingleKey

//SingleKey replaced by SingleKey

//SingleKey replaced by SingleKey

//SingleKey replaced by SingleKey

//SingleKey replaced by SingleKey

//SingleKey replaced by SingleKey

//SingleKey replaced by SingleKey

//SingleKey replaced by SingleKey

//SingleKey replaced by SingleKey

//SingleKey replaced by SingleKey

//SingleKey replaced by SingleKey

//SingleKey replaced by SingleKey

//SingleKey replaced by SingleKey

//SingleKey replaced by SingleKey

//SingleKey replaced by SingleKey

//SingleKey replaced by SingleKey

//SingleKey replaced by SingleKey

//SingleKey replaced by SingleKey

//SingleKey replaced by SingleKey

//SingleKey replaced by SingleKey

//SingleKey replaced by SingleKey

//SingleKey replaced by SingleKey

//SingleKey replaced by SingleKey

//SingleKey replaced by SingleKey

//SingleKey replaced by SingleKey

//SingleKey replaced by SingleKey

//SingleKey replaced by SingleKey

//SingleKey replaced by SingleKey

//SingleKey replaced by SingleKey

//SingleKey replaced by SingleKey

//SingleKey replaced by SingleKey

//SingleKey replaced by SingleKey

//SingleKey replaced by SingleKey

//SingleKey replaced by SingleKey

//SingleKey replaced by SingleKey

//SingleKey replaced by SingleKey

//SingleKey replaced by SingleKey

//SingleKey replaced by SingleKey

//SingleKey replaced by SingleKey

//SingleKey replaced by SingleKey

//SingleKey replaced by SingleKey

//SingleKey replaced by SingleKey

//SingleKey replaced by SingleKey

//SingleKey replaced by SingleKey

//SingleKey replaced by SingleKey

//SingleKey replaced by SingleKey

//SingleKey replaced by SingleKey

//SingleKey replaced by SingleKey

//SingleKey replaced by SingleKey

//SingleKey replaced by SingleKey

//SingleKey replaced by SingleKey

//SingleKey replaced by SingleKey

//SingleKey replaced by SingleKey

//SingleKey replaced by SingleKey

//SingleKey replaced by SingleKey

//SingleKey replaced by SingleKey

//SingleKey replaced by SingleKey

//SingleKey replaced by SingleKey

//SingleKey replaced by SingleKey

//SingleKey replaced by SingleKey

//SingleKey replaced by SingleKey

//SingleKey replaced by SingleKey

//SingleKey replaced by SingleKey

//SingleKey replaced by SingleKey

//SingleKey replaced by SingleKey

//SingleKey replaced by SingleKey

//SingleKey replaced by SingleKey

//SingleKey replaced by SingleKey

//SingleKey replaced by SingleKey

//SingleKey replaced by SingleKey

//SingleKey replaced by SingleKey

//SingleKey replaced by SingleKey

//SingleKey replaced by SingleKey

//SingleKey replaced by SingleKey

//SingleKey replaced by SingleKey

//SingleKey replaced by SingleKey

//SingleKey replaced by SingleKey

//SingleKey replaced by SingleKey

//SingleKey replaced by SingleKey

//SingleKey replaced by SingleKey

//SingleKey replaced by SingleKey

//SingleKey replaced by SingleKey

//SingleKey replaced by SingleKey

//SingleKey replaced by SingleKey

//SingleKey replaced by SingleKey

//SingleKey replaced by SingleKey

//SingleKey replaced by SingleKey

//SingleKey replaced by SingleKey

//SingleKey replaced by SingleKey

//SingleKey replaced by SingleKey

//SingleKey replaced by SingleKey

//SingleKey replaced by SingleKey

//SingleKey replaced by SingleKey

//SingleKey replaced by SingleKey

//SingleKey replaced by SingleKey

module SingleKey (
  input               raw,
  output              filtered_valid,
  output              filtered_payload,
  input               CLK_50,
  input               _zz_3,
  input               _zz_4
);
  reg        [4:0]    cnt;
  reg                 raw_regNext;
  reg                 _zz_1;
  reg                 _zz_2;

  assign filtered_valid = _zz_1;
  assign filtered_payload = _zz_2;
  always @ (posedge CLK_50 or posedge _zz_3) begin
    if (_zz_3) begin
      cnt <= 5'h1a;
    end else begin
      if(_zz_4) begin
        if((raw ^ raw_regNext))begin
          cnt <= 5'h1a;
        end
        if((cnt != 5'h0))begin
          cnt <= (cnt - 5'h01);
        end
      end
    end
  end

  always @ (posedge CLK_50) begin
    if(_zz_4) begin
      raw_regNext <= raw;
      _zz_1 <= (cnt == 5'h01);
      if((cnt == 5'h01))begin
        _zz_2 <= (! raw);
      end
    end
  end


endmodule

module BufferCC (
  input               io_dataIn,
  output              io_dataOut,
  input               CLK_50,
  input               _zz_1
);
  (* async_reg = "true" *) reg                 buffers_0;
  (* async_reg = "true" *) reg                 buffers_1;

  assign io_dataOut = buffers_1;
  always @ (posedge CLK_50 or posedge _zz_1) begin
    if (_zz_1) begin
      buffers_0 <= 1'b0;
      buffers_1 <= 1'b0;
    end else begin
      buffers_0 <= io_dataIn;
      buffers_1 <= buffers_0;
    end
  end


endmodule
