module ps2_rx(
  input clock, clk_in, dat_in, rxen,
  output reg clk_out, dat_out,
  output[7:0] data
);



endmodule
