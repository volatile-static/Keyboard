module ps2_tx(
  input clock, clk_in, dat_in, txen,
  input[7:0] data,
  output reg clk_out, dat_out
);


endmodule
